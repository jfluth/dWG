`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// filename:	icon.v
//
// ECE 540 Project 2: RojoBot World
//
// Jordan Fluth <jfluth@gmail.com>
// Paul Long <pwl@pdx.edu>
//
// 29 October 2014
//
// Description:
//		This module produces the icon that gets painted over the background map
//		produced buy the botsim IP. It relies on the scaling from the 128x128
//		rojobot world to the 512x512 display world to have been done already. 
//		
//		The icon image is stored in a 2D array which is automatically created
//		from an external python script that reads in any bit-mapped image file
//		(.jpg or .png, for example). The array contains the color info for 2 images
//		one pointing North and one pointing NE. The N image is stored in the 256
//		low-order locations and the NE image is stored in the high-order locations.
//		This allows the two Icons to be accessed the same with the exception of the
//		high-order address bit. If that bit is '0', we are addressing the N icon. If 
//		that bit is '1', we are addressing the NE icon.
//		
//		Icons for the other directions are derived on-the-fly by manipulating the
//		order that array is painted onto the screen.
//		
//	General operation:
//		The location reported by the botsim IP is corrected to center the icon
//		on the line. This corrected location is compared to the location of the 
//		cathode ray painting the screen. If the ray is overlapping the bot, the
//		difference between current ray pixel and the bot's top left corner can
//		be used as an index ito the Icon array. The	orientation, as reported by
//		botsim IP, is checked and any necessary	transforms are applied to the
//		indecies to rotate the icon as appropriate.
//
//
//
// 
//
//
//
//////////////////////////////////////////////////////////////////////////////////
module icon (
  
  ///////////////////////////////////////////////////////////////////////////
  // Port Declarations
  ///////////////////////////////////////////////////////////////////////////
  input					clk,
  input			[9:0]	pixCol,			// Current pixel getting drawn
  input			[9:0]	pixRow,
  input			[9:0]	locX,			// RoboCop's current location
  input			[9:0]	locY,			// top left corner
  input			[7:0]	botInfo,
  output	reg	[11:0]	botIcon			// 12-bit rgb color
);


  ///////////////////////////////////////////////////////////////////////////
  // Some Nice Constants
  ///////////////////////////////////////////////////////////////////////////
  localparam N  = 3'b000;				// These are the BotInfo_reg encodings
  localparam S  = 3'b100;				// for compass heading
  localparam E  = 3'b010;
  localparam W  = 3'b110;
  localparam NE = 3'b001;
  localparam SW = 3'b101;
  localparam SE = 3'b011;
  localparam NW = 3'b111;
  //picWidth = 16;
  localparam picwidth = 32;
  
  
  ///////////////////////////////////////////////////////////////////////////
  // Internal Signals
  ///////////////////////////////////////////////////////////////////////////
  reg	[3:0]	iconBitmapX, iconBitmapY;	// index into icon pixelmap 
  wire	[9:0]	iconLeft;					// Bounds of the icon 
  wire	[9:0]	iconRight;
  wire	[9:0]	iconTop;
  wire	[9:0]	iconBottom;
  
  wire	[11:0]	pixelColor;					// Color out from ROM
  reg	[8:0]	romAddress;		
  //reg	[11:0]	iconPixArray[511:0];
  reg [11:0] iconPixArray[2047:0];
 
  
  // These are the icon index transforms that need done in order to use
  // 2 Icons for the eight ordinal directions in which the bot can be headed
  wire	[8:0]	xformN  = {1'b0, 		iconBitmapY,		iconBitmapX }; 
  wire	[8:0]	xformS  = {1'b0, 4'd63-	iconBitmapY, 4'd63-	iconBitmapX }; 
  wire	[8:0]	xformE  = {1'b0, 4'd63-	iconBitmapX, 		iconBitmapY }; 
  wire	[8:0]	xformW  = {1'b0, 		iconBitmapX, 4'd63-	iconBitmapY }; 
  wire	[8:0]	xformNE = {1'b1, 		iconBitmapY, 		iconBitmapX };
  wire	[8:0]	xformSW = {1'b1, 4'd63-	iconBitmapY, 4'd63-	iconBitmapX };
  wire	[8:0]	xformSE = {1'b1, 4'd63-	iconBitmapX, 		iconBitmapY };
  wire	[8:0]	xformNW = {1'b1, 		iconBitmapX, 4'd63-	iconBitmapY };
  
  
  
  ///////////////////////////////////////////////////////////////////////////
  // Global Assigns
  ///////////////////////////////////////////////////////////////////////////
  // This give us an 16x16 box centered on both loc(x,y) and the line
  assign iconLeft   = locX-10'd30; //originl transform is -6 +9
  assign iconRight  = locX+10'd33;
  assign iconTop    = locY-10'd30;
  assign iconBottom = locY+10'd33;
  

  
  // Set index into icon
  always @ (posedge clk) begin
	iconBitmapX <= pixCol[3:0] - iconLeft[3:0];
	iconBitmapY <= pixRow[3:0] -  iconTop[3:0];
  end
  
 
  // Decide when to paint the botIcon
  // If the cathode ray gun overlaps the adjusted bot location,
  // paint the icon, otherwise paint "00" (transparency)

  always @ (posedge clk) begin
	if (pixCol >= iconLeft && pixCol <= iconRight &&
		pixRow >= iconTop  && pixRow <= iconBottom) begin
		
		case (botInfo[2:0])
			N :	botIcon <= iconPixArray[xformN];
			S :	botIcon <= iconPixArray[xformS];
			E :	botIcon <= iconPixArray[xformE];
			W :	botIcon <= iconPixArray[xformW];
			NE:	botIcon <= iconPixArray[xformNE];
			NW:	botIcon <= iconPixArray[xformNW];
			SE:	botIcon <= iconPixArray[xformSE];
			SW:	botIcon <= iconPixArray[xformSW];
			// We should never get here
			default: botIcon <= 12'b0;
		endcase	
	end
	else begin
		botIcon    <= 12'b0;				// transparent 
	end
  end
	  
  initial begin
     /**********************************************
    *****  Template file for the image array
    *****  Produced from icon.png
    ***********************************************/
    iconPixArray[0] = 12'h 00;
    iconPixArray[1] = 12'h 00;
    iconPixArray[2] = 12'h 00;
    iconPixArray[3] = 12'h 00;
    iconPixArray[4] = 12'h 00;
    iconPixArray[5] = 12'h 00;
    iconPixArray[6] = 12'h 00;
    iconPixArray[7] = 12'h247;
    iconPixArray[8] = 12'h246;
    iconPixArray[9] = 12'h 00;
    iconPixArray[10] = 12'h 00;
    iconPixArray[11] = 12'h 00;
    iconPixArray[12] = 12'h 00;
    iconPixArray[13] = 12'h 00;
    iconPixArray[14] = 12'h 00;
    iconPixArray[15] = 12'h 00;
    iconPixArray[16] = 12'h 00;
    iconPixArray[17] = 12'h 00;
    iconPixArray[18] = 12'h 00;
    iconPixArray[19] = 12'h 00;
    iconPixArray[20] = 12'h 00;
    iconPixArray[21] = 12'h 00;
    iconPixArray[22] = 12'h 12;
    iconPixArray[23] = 12'h5AE;
    iconPixArray[24] = 12'h49E;
    iconPixArray[25] = 12'h 11;
    iconPixArray[26] = 12'h 00;
    iconPixArray[27] = 12'h 00;
    iconPixArray[28] = 12'h 00;
    iconPixArray[29] = 12'h 00;
    iconPixArray[30] = 12'h 00;
    iconPixArray[31] = 12'h 00;
    iconPixArray[32] = 12'h 00;
    iconPixArray[33] = 12'h 00;
    iconPixArray[34] = 12'h 00;
    iconPixArray[35] = 12'h 00;
    iconPixArray[36] = 12'h 00;
    iconPixArray[37] = 12'h 00;
    iconPixArray[38] = 12'h36A;
    iconPixArray[39] = 12'h5AF;
    iconPixArray[40] = 12'h5AF;
    iconPixArray[41] = 12'h369;
    iconPixArray[42] = 12'h 00;
    iconPixArray[43] = 12'h 00;
    iconPixArray[44] = 12'h 00;
    iconPixArray[45] = 12'h 00;
    iconPixArray[46] = 12'h 00;
    iconPixArray[47] = 12'h 00;
    iconPixArray[48] = 12'h 00;
    iconPixArray[49] = 12'h 00;
    iconPixArray[50] = 12'h 00;
    iconPixArray[51] = 12'h 00;
    iconPixArray[52] = 12'h 00;
    iconPixArray[53] = 12'h 11;
    iconPixArray[54] = 12'h49E;
    iconPixArray[55] = 12'h49F;
    iconPixArray[56] = 12'h49E;
    iconPixArray[57] = 12'h49E;
    iconPixArray[58] = 12'h 11;
    iconPixArray[59] = 12'h 00;
    iconPixArray[60] = 12'h 00;
    iconPixArray[61] = 12'h 00;
    iconPixArray[62] = 12'h 00;
    iconPixArray[63] = 12'h 00;
    iconPixArray[64] = 12'h 00;
    iconPixArray[65] = 12'h 00;
    iconPixArray[66] = 12'h 00;
    iconPixArray[67] = 12'h 00;
    iconPixArray[68] = 12'h 00;
    iconPixArray[69] = 12'h135;
    iconPixArray[70] = 12'h5AF;
    iconPixArray[71] = 12'h8BE;
    iconPixArray[72] = 12'h9BE;
    iconPixArray[73] = 12'h5AF;
    iconPixArray[74] = 12'h135;
    iconPixArray[75] = 12'h 00;
    iconPixArray[76] = 12'h 00;
    iconPixArray[77] = 12'h 00;
    iconPixArray[78] = 12'h 00;
    iconPixArray[79] = 12'h 00;
    iconPixArray[80] = 12'h 00;
    iconPixArray[81] = 12'h 00;
    iconPixArray[82] = 12'h 00;
    iconPixArray[83] = 12'h 00;
    iconPixArray[84] = 12'h 00;
    iconPixArray[85] = 12'h258;
    iconPixArray[86] = 12'h7BF;
    iconPixArray[87] = 12'hFFE;
    iconPixArray[88] = 12'hFFE;
    iconPixArray[89] = 12'h9CE;
    iconPixArray[90] = 12'h258;
    iconPixArray[91] = 12'h 00;
    iconPixArray[92] = 12'h 00;
    iconPixArray[93] = 12'h 00;
    iconPixArray[94] = 12'h 00;
    iconPixArray[95] = 12'h 00;
    iconPixArray[96] = 12'h 00;
    iconPixArray[97] = 12'h 00;
    iconPixArray[98] = 12'h 00;
    iconPixArray[99] = 12'h 00;
    iconPixArray[100] = 12'h 00;
    iconPixArray[101] = 12'h269;
    iconPixArray[102] = 12'h7BF;
    iconPixArray[103] = 12'hEEE;
    iconPixArray[104] = 12'hFFE;
    iconPixArray[105] = 12'h8CF;
    iconPixArray[106] = 12'h269;
    iconPixArray[107] = 12'h 00;
    iconPixArray[108] = 12'h 00;
    iconPixArray[109] = 12'h 00;
    iconPixArray[110] = 12'h 00;
    iconPixArray[111] = 12'h 00;
    iconPixArray[112] = 12'h 00;
    iconPixArray[113] = 12'h 00;
    iconPixArray[114] = 12'h 00;
    iconPixArray[115] = 12'h 00;
    iconPixArray[116] = 12'h 00;
    iconPixArray[117] = 12'h369;
    iconPixArray[118] = 12'h5AF;
    iconPixArray[119] = 12'h6AE;
    iconPixArray[120] = 12'h7BE;
    iconPixArray[121] = 12'h5AF;
    iconPixArray[122] = 12'h37B;
    iconPixArray[123] = 12'h 00;
    iconPixArray[124] = 12'h 00;
    iconPixArray[125] = 12'h 00;
    iconPixArray[126] = 12'h 00;
    iconPixArray[127] = 12'h 00;
    iconPixArray[128] = 12'h 00;
    iconPixArray[129] = 12'h 00;
    iconPixArray[130] = 12'h 00;
    iconPixArray[131] = 12'h 00;
    iconPixArray[132] = 12'h 00;
    iconPixArray[133] = 12'h269;
    iconPixArray[134] = 12'h5AF;
    iconPixArray[135] = 12'h49E;
    iconPixArray[136] = 12'h49E;
    iconPixArray[137] = 12'h5AF;
    iconPixArray[138] = 12'h26A;
    iconPixArray[139] = 12'h 00;
    iconPixArray[140] = 12'h 00;
    iconPixArray[141] = 12'h 00;
    iconPixArray[142] = 12'h 00;
    iconPixArray[143] = 12'h 00;
    iconPixArray[144] = 12'h 00;
    iconPixArray[145] = 12'h 00;
    iconPixArray[146] = 12'h 00;
    iconPixArray[147] = 12'h 00;
    iconPixArray[148] = 12'h 00;
    iconPixArray[149] = 12'h447;
    iconPixArray[150] = 12'h5AF;
    iconPixArray[151] = 12'h59E;
    iconPixArray[152] = 12'h59E;
    iconPixArray[153] = 12'h4AF;
    iconPixArray[154] = 12'h658;
    iconPixArray[155] = 12'h200;
    iconPixArray[156] = 12'h 00;
    iconPixArray[157] = 12'h 00;
    iconPixArray[158] = 12'h 00;
    iconPixArray[159] = 12'h 00;
    iconPixArray[160] = 12'h 00;
    iconPixArray[161] = 12'h 00;
    iconPixArray[162] = 12'h 00;
    iconPixArray[163] = 12'h 00;
    iconPixArray[164] = 12'h800;
    iconPixArray[165] = 12'hD24;
    iconPixArray[166] = 12'h4AF;
    iconPixArray[167] = 12'h59E;
    iconPixArray[168] = 12'h59E;
    iconPixArray[169] = 12'h4AF;
    iconPixArray[170] = 12'hB47;
    iconPixArray[171] = 12'hD00;
    iconPixArray[172] = 12'h100;
    iconPixArray[173] = 12'h 00;
    iconPixArray[174] = 12'h 00;
    iconPixArray[175] = 12'h 00;
    iconPixArray[176] = 12'h 00;
    iconPixArray[177] = 12'h 00;
    iconPixArray[178] = 12'h 00;
    iconPixArray[179] = 12'h100;
    iconPixArray[180] = 12'hF00;
    iconPixArray[181] = 12'hD12;
    iconPixArray[182] = 12'h59E;
    iconPixArray[183] = 12'h5AF;
    iconPixArray[184] = 12'h59E;
    iconPixArray[185] = 12'h4AE;
    iconPixArray[186] = 12'hB35;
    iconPixArray[187] = 12'hF00;
    iconPixArray[188] = 12'h700;
    iconPixArray[189] = 12'h 00;
    iconPixArray[190] = 12'h 00;
    iconPixArray[191] = 12'h 00;
    iconPixArray[192] = 12'h 00;
    iconPixArray[193] = 12'h 00;
    iconPixArray[194] = 12'h 00;
    iconPixArray[195] = 12'h200;
    iconPixArray[196] = 12'hE00;
    iconPixArray[197] = 12'hE00;
    iconPixArray[198] = 12'h68D;
    iconPixArray[199] = 12'h4AE;
    iconPixArray[200] = 12'h59E;
    iconPixArray[201] = 12'h4AF;
    iconPixArray[202] = 12'hC23;
    iconPixArray[203] = 12'hE00;
    iconPixArray[204] = 12'h600;
    iconPixArray[205] = 12'h 00;
    iconPixArray[206] = 12'h 00;
    iconPixArray[207] = 12'h 00;
    iconPixArray[208] = 12'h 00;
    iconPixArray[209] = 12'h 00;
    iconPixArray[210] = 12'h 00;
    iconPixArray[211] = 12'h 00;
    iconPixArray[212] = 12'hD00;
    iconPixArray[213] = 12'hF00;
    iconPixArray[214] = 12'h78C;
    iconPixArray[215] = 12'h4AF;
    iconPixArray[216] = 12'h59E;
    iconPixArray[217] = 12'h49E;
    iconPixArray[218] = 12'hD12;
    iconPixArray[219] = 12'hF00;
    iconPixArray[220] = 12'h200;
    iconPixArray[221] = 12'h 00;
    iconPixArray[222] = 12'h 00;
    iconPixArray[223] = 12'h 00;
    iconPixArray[224] = 12'h 00;
    iconPixArray[225] = 12'h 00;
    iconPixArray[226] = 12'h 00;
    iconPixArray[227] = 12'h 00;
    iconPixArray[228] = 12'h900;
    iconPixArray[229] = 12'hE00;
    iconPixArray[230] = 12'h223;
    iconPixArray[231] = 12'h123;
    iconPixArray[232] = 12'h112;
    iconPixArray[233] = 12'h 12;
    iconPixArray[234] = 12'h800;
    iconPixArray[235] = 12'hD00;
    iconPixArray[236] = 12'h 00;
    iconPixArray[237] = 12'h 00;
    iconPixArray[238] = 12'h 00;
    iconPixArray[239] = 12'h 00;
    iconPixArray[240] = 12'h 00;
    iconPixArray[241] = 12'h 00;
    iconPixArray[242] = 12'h 00;
    iconPixArray[243] = 12'h 00;
    iconPixArray[244] = 12'h 00;
    iconPixArray[245] = 12'h 00;
    iconPixArray[246] = 12'h 00;
    iconPixArray[247] = 12'h 00;
    iconPixArray[248] = 12'h 00;
    iconPixArray[249] = 12'h 00;
    iconPixArray[250] = 12'h 00;
    iconPixArray[251] = 12'h 00;
    iconPixArray[252] = 12'h 00;
    iconPixArray[253] = 12'h 00;
    iconPixArray[254] = 12'h 00;
    iconPixArray[255] = 12'h 00;
    iconPixArray[256] = 12'h 00;
    iconPixArray[257] = 12'h 00;
    iconPixArray[258] = 12'h 00;
    iconPixArray[259] = 12'h 00;
    iconPixArray[260] = 12'h 00;
    iconPixArray[261] = 12'h 00;
    iconPixArray[262] = 12'h 00;
    iconPixArray[263] = 12'h 00;
    iconPixArray[264] = 12'h 00;
    iconPixArray[265] = 12'h 00;
    iconPixArray[266] = 12'h 00;
    iconPixArray[267] = 12'h 00;
    iconPixArray[268] = 12'h 00;
    iconPixArray[269] = 12'h 00;
    iconPixArray[270] = 12'h 00;
    iconPixArray[271] = 12'h 00;
    iconPixArray[272] = 12'h 00;
    iconPixArray[273] = 12'h 00;
    iconPixArray[274] = 12'h 00;
    iconPixArray[275] = 12'h 00;
    iconPixArray[276] = 12'h 00;
    iconPixArray[277] = 12'h 00;
    iconPixArray[278] = 12'h 00;
    iconPixArray[279] = 12'h 00;
    iconPixArray[280] = 12'h 00;
    iconPixArray[281] = 12'h 00;
    iconPixArray[282] = 12'h 00;
    iconPixArray[283] = 12'h 01;
    iconPixArray[284] = 12'h134;
    iconPixArray[285] = 12'h257;
    iconPixArray[286] = 12'h123;
    iconPixArray[287] = 12'h 00;
    iconPixArray[288] = 12'h 00;
    iconPixArray[289] = 12'h 00;
    iconPixArray[290] = 12'h 00;
    iconPixArray[291] = 12'h 00;
    iconPixArray[292] = 12'h 00;
    iconPixArray[293] = 12'h 00;
    iconPixArray[294] = 12'h 00;
    iconPixArray[295] = 12'h 00;
    iconPixArray[296] = 12'h 00;
    iconPixArray[297] = 12'h 11;
    iconPixArray[298] = 12'h369;
    iconPixArray[299] = 12'h49D;
    iconPixArray[300] = 12'h5AF;
    iconPixArray[301] = 12'h5BF;
    iconPixArray[302] = 12'h124;
    iconPixArray[303] = 12'h 00;
    iconPixArray[304] = 12'h 00;
    iconPixArray[305] = 12'h 00;
    iconPixArray[306] = 12'h 00;
    iconPixArray[307] = 12'h 00;
    iconPixArray[308] = 12'h 00;
    iconPixArray[309] = 12'h 00;
    iconPixArray[310] = 12'h 00;
    iconPixArray[311] = 12'h 00;
    iconPixArray[312] = 12'h135;
    iconPixArray[313] = 12'h49D;
    iconPixArray[314] = 12'h4AF;
    iconPixArray[315] = 12'h49F;
    iconPixArray[316] = 12'h59E;
    iconPixArray[317] = 12'h49E;
    iconPixArray[318] = 12'h 11;
    iconPixArray[319] = 12'h 00;
    iconPixArray[320] = 12'h 00;
    iconPixArray[321] = 12'h 00;
    iconPixArray[322] = 12'h 00;
    iconPixArray[323] = 12'h 00;
    iconPixArray[324] = 12'h 00;
    iconPixArray[325] = 12'h 00;
    iconPixArray[326] = 12'h 00;
    iconPixArray[327] = 12'h246;
    iconPixArray[328] = 12'h5AF;
    iconPixArray[329] = 12'h9CF;
    iconPixArray[330] = 12'hBDE;
    iconPixArray[331] = 12'h7BE;
    iconPixArray[332] = 12'h4AE;
    iconPixArray[333] = 12'h37B;
    iconPixArray[334] = 12'h 00;
    iconPixArray[335] = 12'h 00;
    iconPixArray[336] = 12'h 00;
    iconPixArray[337] = 12'h 00;
    iconPixArray[338] = 12'h 00;
    iconPixArray[339] = 12'h 00;
    iconPixArray[340] = 12'h 00;
    iconPixArray[341] = 12'h 00;
    iconPixArray[342] = 12'h246;
    iconPixArray[343] = 12'h5AF;
    iconPixArray[344] = 12'h5AE;
    iconPixArray[345] = 12'hFEE;
    iconPixArray[346] = 12'hFFF;
    iconPixArray[347] = 12'hCDE;
    iconPixArray[348] = 12'h5AF;
    iconPixArray[349] = 12'h135;
    iconPixArray[350] = 12'h 00;
    iconPixArray[351] = 12'h 00;
    iconPixArray[352] = 12'h 00;
    iconPixArray[353] = 12'h 00;
    iconPixArray[354] = 12'h 00;
    iconPixArray[355] = 12'h600;
    iconPixArray[356] = 12'hA00;
    iconPixArray[357] = 12'h812;
    iconPixArray[358] = 12'h4AE;
    iconPixArray[359] = 12'h5AE;
    iconPixArray[360] = 12'h59E;
    iconPixArray[361] = 12'hBDF;
    iconPixArray[362] = 12'hEEE;
    iconPixArray[363] = 12'h9CF;
    iconPixArray[364] = 12'h37B;
    iconPixArray[365] = 12'h 00;
    iconPixArray[366] = 12'h 00;
    iconPixArray[367] = 12'h 00;
    iconPixArray[368] = 12'h 00;
    iconPixArray[369] = 12'h 00;
    iconPixArray[370] = 12'h600;
    iconPixArray[371] = 12'hF00;
    iconPixArray[372] = 12'hF00;
    iconPixArray[373] = 12'h87B;
    iconPixArray[374] = 12'h4AF;
    iconPixArray[375] = 12'h59E;
    iconPixArray[376] = 12'h49F;
    iconPixArray[377] = 12'h49E;
    iconPixArray[378] = 12'h6AF;
    iconPixArray[379] = 12'h49E;
    iconPixArray[380] = 12'h 11;
    iconPixArray[381] = 12'h 00;
    iconPixArray[382] = 12'h 00;
    iconPixArray[383] = 12'h 00;
    iconPixArray[384] = 12'h 00;
    iconPixArray[385] = 12'h100;
    iconPixArray[386] = 12'hE00;
    iconPixArray[387] = 12'hF00;
    iconPixArray[388] = 12'h957;
    iconPixArray[389] = 12'h4AF;
    iconPixArray[390] = 12'h59E;
    iconPixArray[391] = 12'h5AF;
    iconPixArray[392] = 12'h59E;
    iconPixArray[393] = 12'h5AF;
    iconPixArray[394] = 12'h49E;
    iconPixArray[395] = 12'h123;
    iconPixArray[396] = 12'h 00;
    iconPixArray[397] = 12'h 00;
    iconPixArray[398] = 12'h 00;
    iconPixArray[399] = 12'h 00;
    iconPixArray[400] = 12'h 00;
    iconPixArray[401] = 12'h800;
    iconPixArray[402] = 12'hF00;
    iconPixArray[403] = 12'hC34;
    iconPixArray[404] = 12'h4AE;
    iconPixArray[405] = 12'h59E;
    iconPixArray[406] = 12'h5AE;
    iconPixArray[407] = 12'h59E;
    iconPixArray[408] = 12'h4AF;
    iconPixArray[409] = 12'h49D;
    iconPixArray[410] = 12'h123;
    iconPixArray[411] = 12'h 00;
    iconPixArray[412] = 12'h 00;
    iconPixArray[413] = 12'h 00;
    iconPixArray[414] = 12'h 00;
    iconPixArray[415] = 12'h 00;
    iconPixArray[416] = 12'h 00;
    iconPixArray[417] = 12'h700;
    iconPixArray[418] = 12'h400;
    iconPixArray[419] = 12'h258;
    iconPixArray[420] = 12'h5AF;
    iconPixArray[421] = 12'h59E;
    iconPixArray[422] = 12'h59E;
    iconPixArray[423] = 12'h4AF;
    iconPixArray[424] = 12'h87B;
    iconPixArray[425] = 12'hB11;
    iconPixArray[426] = 12'h 00;
    iconPixArray[427] = 12'h 00;
    iconPixArray[428] = 12'h 00;
    iconPixArray[429] = 12'h 00;
    iconPixArray[430] = 12'h 00;
    iconPixArray[431] = 12'h 00;
    iconPixArray[432] = 12'h 00;
    iconPixArray[433] = 12'h 00;
    iconPixArray[434] = 12'h 00;
    iconPixArray[435] = 12'h 00;
    iconPixArray[436] = 12'h258;
    iconPixArray[437] = 12'h5AF;
    iconPixArray[438] = 12'h4AF;
    iconPixArray[439] = 12'h958;
    iconPixArray[440] = 12'hE00;
    iconPixArray[441] = 12'hD00;
    iconPixArray[442] = 12'h 00;
    iconPixArray[443] = 12'h 00;
    iconPixArray[444] = 12'h 00;
    iconPixArray[445] = 12'h 00;
    iconPixArray[446] = 12'h 00;
    iconPixArray[447] = 12'h 00;
    iconPixArray[448] = 12'h 00;
    iconPixArray[449] = 12'h 00;
    iconPixArray[450] = 12'h 00;
    iconPixArray[451] = 12'h 00;
    iconPixArray[452] = 12'h 00;
    iconPixArray[453] = 12'h157;
    iconPixArray[454] = 12'hA46;
    iconPixArray[455] = 12'hF00;
    iconPixArray[456] = 12'hF00;
    iconPixArray[457] = 12'h800;
    iconPixArray[458] = 12'h 00;
    iconPixArray[459] = 12'h 00;
    iconPixArray[460] = 12'h 00;
    iconPixArray[461] = 12'h 00;
    iconPixArray[462] = 12'h 00;
    iconPixArray[463] = 12'h 00;
    iconPixArray[464] = 12'h 00;
    iconPixArray[465] = 12'h 00;
    iconPixArray[466] = 12'h 00;
    iconPixArray[467] = 12'h 00;
    iconPixArray[468] = 12'h 00;
    iconPixArray[469] = 12'h100;
    iconPixArray[470] = 12'hF00;
    iconPixArray[471] = 12'hE00;
    iconPixArray[472] = 12'h800;
    iconPixArray[473] = 12'h 00;
    iconPixArray[474] = 12'h 00;
    iconPixArray[475] = 12'h 00;
    iconPixArray[476] = 12'h 00;
    iconPixArray[477] = 12'h 00;
    iconPixArray[478] = 12'h 00;
    iconPixArray[479] = 12'h 00;
    iconPixArray[480] = 12'h 00;
    iconPixArray[481] = 12'h 00;
    iconPixArray[482] = 12'h 00;
    iconPixArray[483] = 12'h 00;
    iconPixArray[484] = 12'h 00;
    iconPixArray[485] = 12'h400;
    iconPixArray[486] = 12'h800;
    iconPixArray[487] = 12'h200;
    iconPixArray[488] = 12'h 00;
    iconPixArray[489] = 12'h 00;
    iconPixArray[490] = 12'h 00;
    iconPixArray[491] = 12'h 00;
    iconPixArray[492] = 12'h 00;
    iconPixArray[493] = 12'h 00;
    iconPixArray[494] = 12'h 00;
    iconPixArray[495] = 12'h 00;
    iconPixArray[496] = 12'h 00;
    iconPixArray[497] = 12'h 00;
    iconPixArray[498] = 12'h 00;
    iconPixArray[499] = 12'h 00;
    iconPixArray[500] = 12'h 00;
    iconPixArray[501] = 12'h 00;
    iconPixArray[502] = 12'h 00;
    iconPixArray[503] = 12'h 00;
    iconPixArray[504] = 12'h 00;
    iconPixArray[505] = 12'h 00;
    iconPixArray[506] = 12'h 00;
    iconPixArray[507] = 12'h 00;
    iconPixArray[508] = 12'h 00;
    iconPixArray[509] = 12'h 00;
    iconPixArray[510] = 12'h 00;
    iconPixArray[511] = 12'h 00;

/**********************************************
*****  Template file for the image array
*****  Produced from fireRocket.png
***********************************************/
/*
iconPixArray[0] = 12'h 00;
iconPixArray[1] = 12'h 00;
iconPixArray[2] = 12'h 00;
iconPixArray[3] = 12'h 00;
iconPixArray[4] = 12'h 00;
iconPixArray[5] = 12'h 00;
iconPixArray[6] = 12'h 00;
iconPixArray[7] = 12'h 00;
iconPixArray[8] = 12'h 00;
iconPixArray[9] = 12'h 00;
iconPixArray[10] = 12'h 00;
iconPixArray[11] = 12'h 00;
iconPixArray[12] = 12'h 00;
iconPixArray[13] = 12'h 00;
iconPixArray[14] = 12'h 00;
iconPixArray[15] = 12'h 00;
iconPixArray[16] = 12'h 00;
iconPixArray[17] = 12'h 00;
iconPixArray[18] = 12'h 00;
iconPixArray[19] = 12'h 00;
iconPixArray[20] = 12'h 00;
iconPixArray[21] = 12'h 00;
iconPixArray[22] = 12'h 00;
iconPixArray[23] = 12'h 00;
iconPixArray[24] = 12'h 00;
iconPixArray[25] = 12'h 00;
iconPixArray[26] = 12'h 00;
iconPixArray[27] = 12'h 00;
iconPixArray[28] = 12'h 00;
iconPixArray[29] = 12'h 00;
iconPixArray[30] = 12'h 00;
iconPixArray[31] = 12'h 00;
iconPixArray[32] = 12'h 00;
iconPixArray[33] = 12'h 00;
iconPixArray[34] = 12'h 00;
iconPixArray[35] = 12'h 00;
iconPixArray[36] = 12'h 00;
iconPixArray[37] = 12'h 00;
iconPixArray[38] = 12'h 00;
iconPixArray[39] = 12'h 00;
iconPixArray[40] = 12'h 00;
iconPixArray[41] = 12'h 00;
iconPixArray[42] = 12'h 00;
iconPixArray[43] = 12'h 00;
iconPixArray[44] = 12'h 00;
iconPixArray[45] = 12'h 00;
iconPixArray[46] = 12'h 00;
iconPixArray[47] = 12'h 00;
iconPixArray[48] = 12'h 00;
iconPixArray[49] = 12'h 00;
iconPixArray[50] = 12'h 00;
iconPixArray[51] = 12'h 00;
iconPixArray[52] = 12'h 00;
iconPixArray[53] = 12'h 00;
iconPixArray[54] = 12'h 00;
iconPixArray[55] = 12'h 00;
iconPixArray[56] = 12'h 00;
iconPixArray[57] = 12'h 00;
iconPixArray[58] = 12'h 00;
iconPixArray[59] = 12'h 00;
iconPixArray[60] = 12'h 00;
iconPixArray[61] = 12'h 00;
iconPixArray[62] = 12'h 00;
iconPixArray[63] = 12'h 00;
iconPixArray[64] = 12'h 00;
iconPixArray[65] = 12'h 00;
iconPixArray[66] = 12'h 00;
iconPixArray[67] = 12'h 00;
iconPixArray[68] = 12'h 00;
iconPixArray[69] = 12'h 00;
iconPixArray[70] = 12'h 00;
iconPixArray[71] = 12'h 00;
iconPixArray[72] = 12'h 00;
iconPixArray[73] = 12'h 00;
iconPixArray[74] = 12'h 00;
iconPixArray[75] = 12'h 00;
iconPixArray[76] = 12'h 00;
iconPixArray[77] = 12'h 00;
iconPixArray[78] = 12'h 00;
iconPixArray[79] = 12'h333;
iconPixArray[80] = 12'h999;
iconPixArray[81] = 12'h 00;
iconPixArray[82] = 12'h 00;
iconPixArray[83] = 12'h 00;
iconPixArray[84] = 12'h 00;
iconPixArray[85] = 12'h 00;
iconPixArray[86] = 12'h 00;
iconPixArray[87] = 12'h 00;
iconPixArray[88] = 12'h 00;
iconPixArray[89] = 12'h 00;
iconPixArray[90] = 12'h 00;
iconPixArray[91] = 12'h 00;
iconPixArray[92] = 12'h 00;
iconPixArray[93] = 12'h 00;
iconPixArray[94] = 12'h 00;
iconPixArray[95] = 12'h 00;
iconPixArray[96] = 12'h 00;
iconPixArray[97] = 12'h 00;
iconPixArray[98] = 12'h 00;
iconPixArray[99] = 12'h 00;
iconPixArray[100] = 12'h 00;
iconPixArray[101] = 12'h 00;
iconPixArray[102] = 12'h 00;
iconPixArray[103] = 12'h 00;
iconPixArray[104] = 12'h 00;
iconPixArray[105] = 12'h 00;
iconPixArray[106] = 12'h 00;
iconPixArray[107] = 12'h 00;
iconPixArray[108] = 12'h 00;
iconPixArray[109] = 12'h 00;
iconPixArray[110] = 12'h 00;
iconPixArray[111] = 12'hBBB;
iconPixArray[112] = 12'hEEE;
iconPixArray[113] = 12'h666;
iconPixArray[114] = 12'h 00;
iconPixArray[115] = 12'h 00;
iconPixArray[116] = 12'h 00;
iconPixArray[117] = 12'h 00;
iconPixArray[118] = 12'h 00;
iconPixArray[119] = 12'h 00;
iconPixArray[120] = 12'h 00;
iconPixArray[121] = 12'h 00;
iconPixArray[122] = 12'h 00;
iconPixArray[123] = 12'h 00;
iconPixArray[124] = 12'h 00;
iconPixArray[125] = 12'h 00;
iconPixArray[126] = 12'h 00;
iconPixArray[127] = 12'h 00;
iconPixArray[128] = 12'h 00;
iconPixArray[129] = 12'h 00;
iconPixArray[130] = 12'h 00;
iconPixArray[131] = 12'h 00;
iconPixArray[132] = 12'h 00;
iconPixArray[133] = 12'h 00;
iconPixArray[134] = 12'h 00;
iconPixArray[135] = 12'h 00;
iconPixArray[136] = 12'h 00;
iconPixArray[137] = 12'h 00;
iconPixArray[138] = 12'h 00;
iconPixArray[139] = 12'h 00;
iconPixArray[140] = 12'h 00;
iconPixArray[141] = 12'h 00;
iconPixArray[142] = 12'h666;
iconPixArray[143] = 12'hDDD;
iconPixArray[144] = 12'hCCC;
iconPixArray[145] = 12'hCCC;
iconPixArray[146] = 12'h222;
iconPixArray[147] = 12'h 00;
iconPixArray[148] = 12'h 00;
iconPixArray[149] = 12'h 00;
iconPixArray[150] = 12'h 00;
iconPixArray[151] = 12'h 00;
iconPixArray[152] = 12'h 00;
iconPixArray[153] = 12'h 00;
iconPixArray[154] = 12'h 00;
iconPixArray[155] = 12'h 00;
iconPixArray[156] = 12'h 00;
iconPixArray[157] = 12'h 00;
iconPixArray[158] = 12'h 00;
iconPixArray[159] = 12'h 00;
iconPixArray[160] = 12'h 00;
iconPixArray[161] = 12'h 00;
iconPixArray[162] = 12'h 00;
iconPixArray[163] = 12'h 00;
iconPixArray[164] = 12'h 00;
iconPixArray[165] = 12'h 00;
iconPixArray[166] = 12'h 00;
iconPixArray[167] = 12'h 00;
iconPixArray[168] = 12'h 00;
iconPixArray[169] = 12'h 00;
iconPixArray[170] = 12'h 00;
iconPixArray[171] = 12'h 00;
iconPixArray[172] = 12'h 00;
iconPixArray[173] = 12'h111;
iconPixArray[174] = 12'hCCC;
iconPixArray[175] = 12'hCCC;
iconPixArray[176] = 12'hCCC;
iconPixArray[177] = 12'hDDD;
iconPixArray[178] = 12'h888;
iconPixArray[179] = 12'h 00;
iconPixArray[180] = 12'h 00;
iconPixArray[181] = 12'h 00;
iconPixArray[182] = 12'h 00;
iconPixArray[183] = 12'h 00;
iconPixArray[184] = 12'h 00;
iconPixArray[185] = 12'h 00;
iconPixArray[186] = 12'h 00;
iconPixArray[187] = 12'h 00;
iconPixArray[188] = 12'h 00;
iconPixArray[189] = 12'h 00;
iconPixArray[190] = 12'h 00;
iconPixArray[191] = 12'h 00;
iconPixArray[192] = 12'h 00;
iconPixArray[193] = 12'h 00;
iconPixArray[194] = 12'h 00;
iconPixArray[195] = 12'h 00;
iconPixArray[196] = 12'h 00;
iconPixArray[197] = 12'h 00;
iconPixArray[198] = 12'h 00;
iconPixArray[199] = 12'h 00;
iconPixArray[200] = 12'h 00;
iconPixArray[201] = 12'h 00;
iconPixArray[202] = 12'h 00;
iconPixArray[203] = 12'h 00;
iconPixArray[204] = 12'h 00;
iconPixArray[205] = 12'h666;
iconPixArray[206] = 12'hDDD;
iconPixArray[207] = 12'hCCC;
iconPixArray[208] = 12'hDDD;
iconPixArray[209] = 12'hCCC;
iconPixArray[210] = 12'hDDD;
iconPixArray[211] = 12'h222;
iconPixArray[212] = 12'h 00;
iconPixArray[213] = 12'h 00;
iconPixArray[214] = 12'h 00;
iconPixArray[215] = 12'h 00;
iconPixArray[216] = 12'h 00;
iconPixArray[217] = 12'h 00;
iconPixArray[218] = 12'h 00;
iconPixArray[219] = 12'h 00;
iconPixArray[220] = 12'h 00;
iconPixArray[221] = 12'h 00;
iconPixArray[222] = 12'h 00;
iconPixArray[223] = 12'h 00;
iconPixArray[224] = 12'h 00;
iconPixArray[225] = 12'h 00;
iconPixArray[226] = 12'h 00;
iconPixArray[227] = 12'h 00;
iconPixArray[228] = 12'h 00;
iconPixArray[229] = 12'h 00;
iconPixArray[230] = 12'h 00;
iconPixArray[231] = 12'h 00;
iconPixArray[232] = 12'h 00;
iconPixArray[233] = 12'h 00;
iconPixArray[234] = 12'h 00;
iconPixArray[235] = 12'h 00;
iconPixArray[236] = 12'h 00;
iconPixArray[237] = 12'hAAA;
iconPixArray[238] = 12'hDDD;
iconPixArray[239] = 12'hCCC;
iconPixArray[240] = 12'hBBB;
iconPixArray[241] = 12'hDDD;
iconPixArray[242] = 12'hDDD;
iconPixArray[243] = 12'h777;
iconPixArray[244] = 12'h 00;
iconPixArray[245] = 12'h 00;
iconPixArray[246] = 12'h 00;
iconPixArray[247] = 12'h 00;
iconPixArray[248] = 12'h 00;
iconPixArray[249] = 12'h 00;
iconPixArray[250] = 12'h 00;
iconPixArray[251] = 12'h 00;
iconPixArray[252] = 12'h 00;
iconPixArray[253] = 12'h 00;
iconPixArray[254] = 12'h 00;
iconPixArray[255] = 12'h 00;
iconPixArray[256] = 12'h 00;
iconPixArray[257] = 12'h 00;
iconPixArray[258] = 12'h 00;
iconPixArray[259] = 12'h 00;
iconPixArray[260] = 12'h 00;
iconPixArray[261] = 12'h 00;
iconPixArray[262] = 12'h 00;
iconPixArray[263] = 12'h 00;
iconPixArray[264] = 12'h 00;
iconPixArray[265] = 12'h 00;
iconPixArray[266] = 12'h 00;
iconPixArray[267] = 12'h 00;
iconPixArray[268] = 12'h222;
iconPixArray[269] = 12'hDDD;
iconPixArray[270] = 12'hAAA;
iconPixArray[271] = 12'h222;
iconPixArray[272] = 12'h222;
iconPixArray[273] = 12'h666;
iconPixArray[274] = 12'hDDD;
iconPixArray[275] = 12'hBBB;
iconPixArray[276] = 12'h 00;
iconPixArray[277] = 12'h 00;
iconPixArray[278] = 12'h 00;
iconPixArray[279] = 12'h 00;
iconPixArray[280] = 12'h 00;
iconPixArray[281] = 12'h 00;
iconPixArray[282] = 12'h 00;
iconPixArray[283] = 12'h 00;
iconPixArray[284] = 12'h 00;
iconPixArray[285] = 12'h 00;
iconPixArray[286] = 12'h 00;
iconPixArray[287] = 12'h 00;
iconPixArray[288] = 12'h 00;
iconPixArray[289] = 12'h 00;
iconPixArray[290] = 12'h 00;
iconPixArray[291] = 12'h 00;
iconPixArray[292] = 12'h 00;
iconPixArray[293] = 12'h 00;
iconPixArray[294] = 12'h 00;
iconPixArray[295] = 12'h 00;
iconPixArray[296] = 12'h 00;
iconPixArray[297] = 12'h 00;
iconPixArray[298] = 12'h 00;
iconPixArray[299] = 12'h 00;
iconPixArray[300] = 12'h444;
iconPixArray[301] = 12'hEEE;
iconPixArray[302] = 12'h444;
iconPixArray[303] = 12'h799;
iconPixArray[304] = 12'hBDD;
iconPixArray[305] = 12'h222;
iconPixArray[306] = 12'hAAA;
iconPixArray[307] = 12'hDDD;
iconPixArray[308] = 12'h333;
iconPixArray[309] = 12'h 00;
iconPixArray[310] = 12'h 00;
iconPixArray[311] = 12'h 00;
iconPixArray[312] = 12'h 00;
iconPixArray[313] = 12'h 00;
iconPixArray[314] = 12'h 00;
iconPixArray[315] = 12'h 00;
iconPixArray[316] = 12'h 00;
iconPixArray[317] = 12'h 00;
iconPixArray[318] = 12'h 00;
iconPixArray[319] = 12'h 00;
iconPixArray[320] = 12'h 00;
iconPixArray[321] = 12'h 00;
iconPixArray[322] = 12'h 00;
iconPixArray[323] = 12'h 00;
iconPixArray[324] = 12'h 00;
iconPixArray[325] = 12'h 00;
iconPixArray[326] = 12'h 00;
iconPixArray[327] = 12'h 00;
iconPixArray[328] = 12'h 00;
iconPixArray[329] = 12'h 00;
iconPixArray[330] = 12'h 00;
iconPixArray[331] = 12'h 00;
iconPixArray[332] = 12'h777;
iconPixArray[333] = 12'hEEE;
iconPixArray[334] = 12'h444;
iconPixArray[335] = 12'h688;
iconPixArray[336] = 12'hBDD;
iconPixArray[337] = 12'h222;
iconPixArray[338] = 12'hAAA;
iconPixArray[339] = 12'hEEE;
iconPixArray[340] = 12'h666;
iconPixArray[341] = 12'h 00;
iconPixArray[342] = 12'h 00;
iconPixArray[343] = 12'h 00;
iconPixArray[344] = 12'h 00;
iconPixArray[345] = 12'h 00;
iconPixArray[346] = 12'h 00;
iconPixArray[347] = 12'h 00;
iconPixArray[348] = 12'h 00;
iconPixArray[349] = 12'h 00;
iconPixArray[350] = 12'h 00;
iconPixArray[351] = 12'h 00;
iconPixArray[352] = 12'h 00;
iconPixArray[353] = 12'h 00;
iconPixArray[354] = 12'h 00;
iconPixArray[355] = 12'h 00;
iconPixArray[356] = 12'h 00;
iconPixArray[357] = 12'h 00;
iconPixArray[358] = 12'h 00;
iconPixArray[359] = 12'h 00;
iconPixArray[360] = 12'h 00;
iconPixArray[361] = 12'h 00;
iconPixArray[362] = 12'h 00;
iconPixArray[363] = 12'h 00;
iconPixArray[364] = 12'h888;
iconPixArray[365] = 12'hEEE;
iconPixArray[366] = 12'hAAA;
iconPixArray[367] = 12'h222;
iconPixArray[368] = 12'h222;
iconPixArray[369] = 12'h666;
iconPixArray[370] = 12'hDDD;
iconPixArray[371] = 12'hDDD;
iconPixArray[372] = 12'h888;
iconPixArray[373] = 12'h 00;
iconPixArray[374] = 12'h 00;
iconPixArray[375] = 12'h 00;
iconPixArray[376] = 12'h 00;
iconPixArray[377] = 12'h 00;
iconPixArray[378] = 12'h 00;
iconPixArray[379] = 12'h 00;
iconPixArray[380] = 12'h 00;
iconPixArray[381] = 12'h 00;
iconPixArray[382] = 12'h 00;
iconPixArray[383] = 12'h 00;
iconPixArray[384] = 12'h 00;
iconPixArray[385] = 12'h 00;
iconPixArray[386] = 12'h 00;
iconPixArray[387] = 12'h 00;
iconPixArray[388] = 12'h 00;
iconPixArray[389] = 12'h 00;
iconPixArray[390] = 12'h 00;
iconPixArray[391] = 12'h 00;
iconPixArray[392] = 12'h 00;
iconPixArray[393] = 12'h 00;
iconPixArray[394] = 12'h 00;
iconPixArray[395] = 12'h 00;
iconPixArray[396] = 12'h999;
iconPixArray[397] = 12'hDDD;
iconPixArray[398] = 12'hDDD;
iconPixArray[399] = 12'hCCC;
iconPixArray[400] = 12'hBBB;
iconPixArray[401] = 12'hDDD;
iconPixArray[402] = 12'hCCC;
iconPixArray[403] = 12'hDDD;
iconPixArray[404] = 12'h999;
iconPixArray[405] = 12'h 00;
iconPixArray[406] = 12'h 00;
iconPixArray[407] = 12'h 00;
iconPixArray[408] = 12'h 00;
iconPixArray[409] = 12'h 00;
iconPixArray[410] = 12'h 00;
iconPixArray[411] = 12'h 00;
iconPixArray[412] = 12'h 00;
iconPixArray[413] = 12'h 00;
iconPixArray[414] = 12'h 00;
iconPixArray[415] = 12'h 00;
iconPixArray[416] = 12'h 00;
iconPixArray[417] = 12'h 00;
iconPixArray[418] = 12'h 00;
iconPixArray[419] = 12'h 00;
iconPixArray[420] = 12'h 00;
iconPixArray[421] = 12'h 00;
iconPixArray[422] = 12'h 00;
iconPixArray[423] = 12'h 00;
iconPixArray[424] = 12'h 00;
iconPixArray[425] = 12'h 00;
iconPixArray[426] = 12'h 00;
iconPixArray[427] = 12'h 00;
iconPixArray[428] = 12'hAAA;
iconPixArray[429] = 12'hDDD;
iconPixArray[430] = 12'hCCC;
iconPixArray[431] = 12'hCCC;
iconPixArray[432] = 12'hCCC;
iconPixArray[433] = 12'hCCC;
iconPixArray[434] = 12'hCCC;
iconPixArray[435] = 12'hDDD;
iconPixArray[436] = 12'h999;
iconPixArray[437] = 12'h 00;
iconPixArray[438] = 12'h 00;
iconPixArray[439] = 12'h 00;
iconPixArray[440] = 12'h 00;
iconPixArray[441] = 12'h 00;
iconPixArray[442] = 12'h 00;
iconPixArray[443] = 12'h 00;
iconPixArray[444] = 12'h 00;
iconPixArray[445] = 12'h 00;
iconPixArray[446] = 12'h 00;
iconPixArray[447] = 12'h 00;
iconPixArray[448] = 12'h 00;
iconPixArray[449] = 12'h 00;
iconPixArray[450] = 12'h 00;
iconPixArray[451] = 12'h 00;
iconPixArray[452] = 12'h 00;
iconPixArray[453] = 12'h 00;
iconPixArray[454] = 12'h 00;
iconPixArray[455] = 12'h 00;
iconPixArray[456] = 12'h 00;
iconPixArray[457] = 12'h 00;
iconPixArray[458] = 12'h 00;
iconPixArray[459] = 12'h 00;
iconPixArray[460] = 12'hAAA;
iconPixArray[461] = 12'hDDD;
iconPixArray[462] = 12'hCCC;
iconPixArray[463] = 12'h666;
iconPixArray[464] = 12'h333;
iconPixArray[465] = 12'hAAA;
iconPixArray[466] = 12'hDDD;
iconPixArray[467] = 12'hDDD;
iconPixArray[468] = 12'h999;
iconPixArray[469] = 12'h 00;
iconPixArray[470] = 12'h 00;
iconPixArray[471] = 12'h 00;
iconPixArray[472] = 12'h 00;
iconPixArray[473] = 12'h 00;
iconPixArray[474] = 12'h 00;
iconPixArray[475] = 12'h 00;
iconPixArray[476] = 12'h 00;
iconPixArray[477] = 12'h 00;
iconPixArray[478] = 12'h 00;
iconPixArray[479] = 12'h 00;
iconPixArray[480] = 12'h 00;
iconPixArray[481] = 12'h 00;
iconPixArray[482] = 12'h 00;
iconPixArray[483] = 12'h 00;
iconPixArray[484] = 12'h 00;
iconPixArray[485] = 12'h 00;
iconPixArray[486] = 12'h 00;
iconPixArray[487] = 12'h 00;
iconPixArray[488] = 12'h 00;
iconPixArray[489] = 12'h 00;
iconPixArray[490] = 12'h111;
iconPixArray[491] = 12'h555;
iconPixArray[492] = 12'h999;
iconPixArray[493] = 12'hEEE;
iconPixArray[494] = 12'hAAA;
iconPixArray[495] = 12'h666;
iconPixArray[496] = 12'h333;
iconPixArray[497] = 12'hAAA;
iconPixArray[498] = 12'hDDD;
iconPixArray[499] = 12'hDDD;
iconPixArray[500] = 12'h888;
iconPixArray[501] = 12'h111;
iconPixArray[502] = 12'h 00;
iconPixArray[503] = 12'h 00;
iconPixArray[504] = 12'h 00;
iconPixArray[505] = 12'h 00;
iconPixArray[506] = 12'h 00;
iconPixArray[507] = 12'h 00;
iconPixArray[508] = 12'h 00;
iconPixArray[509] = 12'h 00;
iconPixArray[510] = 12'h 00;
iconPixArray[511] = 12'h 00;
iconPixArray[512] = 12'h 00;
iconPixArray[513] = 12'h 00;
iconPixArray[514] = 12'h 00;
iconPixArray[515] = 12'h 00;
iconPixArray[516] = 12'h 00;
iconPixArray[517] = 12'h 00;
iconPixArray[518] = 12'h 00;
iconPixArray[519] = 12'h 00;
iconPixArray[520] = 12'h 00;
iconPixArray[521] = 12'h111;
iconPixArray[522] = 12'h999;
iconPixArray[523] = 12'h999;
iconPixArray[524] = 12'h888;
iconPixArray[525] = 12'hEEE;
iconPixArray[526] = 12'h999;
iconPixArray[527] = 12'h666;
iconPixArray[528] = 12'h444;
iconPixArray[529] = 12'hAAA;
iconPixArray[530] = 12'hDDD;
iconPixArray[531] = 12'hDDD;
iconPixArray[532] = 12'h777;
iconPixArray[533] = 12'h999;
iconPixArray[534] = 12'h111;
iconPixArray[535] = 12'h 00;
iconPixArray[536] = 12'h 00;
iconPixArray[537] = 12'h 00;
iconPixArray[538] = 12'h 00;
iconPixArray[539] = 12'h 00;
iconPixArray[540] = 12'h 00;
iconPixArray[541] = 12'h 00;
iconPixArray[542] = 12'h 00;
iconPixArray[543] = 12'h 00;
iconPixArray[544] = 12'h 00;
iconPixArray[545] = 12'h 00;
iconPixArray[546] = 12'h 00;
iconPixArray[547] = 12'h 00;
iconPixArray[548] = 12'h 00;
iconPixArray[549] = 12'h 00;
iconPixArray[550] = 12'h 00;
iconPixArray[551] = 12'h 00;
iconPixArray[552] = 12'h 00;
iconPixArray[553] = 12'h555;
iconPixArray[554] = 12'hCCC;
iconPixArray[555] = 12'h999;
iconPixArray[556] = 12'h777;
iconPixArray[557] = 12'hDDD;
iconPixArray[558] = 12'h999;
iconPixArray[559] = 12'h666;
iconPixArray[560] = 12'h444;
iconPixArray[561] = 12'hAAA;
iconPixArray[562] = 12'hDDD;
iconPixArray[563] = 12'hCCC;
iconPixArray[564] = 12'h666;
iconPixArray[565] = 12'hBBB;
iconPixArray[566] = 12'h999;
iconPixArray[567] = 12'h 00;
iconPixArray[568] = 12'h 00;
iconPixArray[569] = 12'h 00;
iconPixArray[570] = 12'h 00;
iconPixArray[571] = 12'h 00;
iconPixArray[572] = 12'h 00;
iconPixArray[573] = 12'h 00;
iconPixArray[574] = 12'h 00;
iconPixArray[575] = 12'h 00;
iconPixArray[576] = 12'h 00;
iconPixArray[577] = 12'h 00;
iconPixArray[578] = 12'h 00;
iconPixArray[579] = 12'h 00;
iconPixArray[580] = 12'h 00;
iconPixArray[581] = 12'h 00;
iconPixArray[582] = 12'h 00;
iconPixArray[583] = 12'h 00;
iconPixArray[584] = 12'h 00;
iconPixArray[585] = 12'h222;
iconPixArray[586] = 12'hBBB;
iconPixArray[587] = 12'hAAA;
iconPixArray[588] = 12'h666;
iconPixArray[589] = 12'hEEE;
iconPixArray[590] = 12'hAAB;
iconPixArray[591] = 12'h666;
iconPixArray[592] = 12'h444;
iconPixArray[593] = 12'hBBB;
iconPixArray[594] = 12'hEEE;
iconPixArray[595] = 12'hAAA;
iconPixArray[596] = 12'h666;
iconPixArray[597] = 12'hCCC;
iconPixArray[598] = 12'hAAA;
iconPixArray[599] = 12'h 00;
iconPixArray[600] = 12'h 00;
iconPixArray[601] = 12'h 00;
iconPixArray[602] = 12'h 00;
iconPixArray[603] = 12'h 00;
iconPixArray[604] = 12'h 00;
iconPixArray[605] = 12'h 00;
iconPixArray[606] = 12'h 00;
iconPixArray[607] = 12'h 00;
iconPixArray[608] = 12'h 00;
iconPixArray[609] = 12'h 00;
iconPixArray[610] = 12'h 00;
iconPixArray[611] = 12'h 00;
iconPixArray[612] = 12'h 00;
iconPixArray[613] = 12'h 00;
iconPixArray[614] = 12'h 00;
iconPixArray[615] = 12'h 00;
iconPixArray[616] = 12'h 00;
iconPixArray[617] = 12'h 00;
iconPixArray[618] = 12'h999;
iconPixArray[619] = 12'hCCC;
iconPixArray[620] = 12'h666;
iconPixArray[621] = 12'h888;
iconPixArray[622] = 12'h666;
iconPixArray[623] = 12'h666;
iconPixArray[624] = 12'h344;
iconPixArray[625] = 12'h666;
iconPixArray[626] = 12'hABB;
iconPixArray[627] = 12'h677;
iconPixArray[628] = 12'h999;
iconPixArray[629] = 12'hCCC;
iconPixArray[630] = 12'h555;
iconPixArray[631] = 12'h 00;
iconPixArray[632] = 12'h 00;
iconPixArray[633] = 12'h 00;
iconPixArray[634] = 12'h 00;
iconPixArray[635] = 12'h 00;
iconPixArray[636] = 12'h 00;
iconPixArray[637] = 12'h 00;
iconPixArray[638] = 12'h 00;
iconPixArray[639] = 12'h 00;
iconPixArray[640] = 12'h 00;
iconPixArray[641] = 12'h 00;
iconPixArray[642] = 12'h 00;
iconPixArray[643] = 12'h 00;
iconPixArray[644] = 12'h 00;
iconPixArray[645] = 12'h 00;
iconPixArray[646] = 12'h 00;
iconPixArray[647] = 12'h 00;
iconPixArray[648] = 12'h 00;
iconPixArray[649] = 12'h 00;
iconPixArray[650] = 12'h777;
iconPixArray[651] = 12'hBCC;
iconPixArray[652] = 12'h522;
iconPixArray[653] = 12'hB50;
iconPixArray[654] = 12'hB90;
iconPixArray[655] = 12'h444;
iconPixArray[656] = 12'h432;
iconPixArray[657] = 12'hB91;
iconPixArray[658] = 12'h930;
iconPixArray[659] = 12'h422;
iconPixArray[660] = 12'hBBB;
iconPixArray[661] = 12'hAAA;
iconPixArray[662] = 12'h111;
iconPixArray[663] = 12'h 00;
iconPixArray[664] = 12'h 00;
iconPixArray[665] = 12'h 00;
iconPixArray[666] = 12'h 00;
iconPixArray[667] = 12'h 00;
iconPixArray[668] = 12'h 00;
iconPixArray[669] = 12'h 00;
iconPixArray[670] = 12'h 00;
iconPixArray[671] = 12'h 00;
iconPixArray[672] = 12'h 00;
iconPixArray[673] = 12'h 00;
iconPixArray[674] = 12'h 00;
iconPixArray[675] = 12'h 00;
iconPixArray[676] = 12'h 00;
iconPixArray[677] = 12'h 00;
iconPixArray[678] = 12'h 00;
iconPixArray[679] = 12'h 00;
iconPixArray[680] = 12'h 00;
iconPixArray[681] = 12'h 00;
iconPixArray[682] = 12'h333;
iconPixArray[683] = 12'h434;
iconPixArray[684] = 12'hB30;
iconPixArray[685] = 12'hFC2;
iconPixArray[686] = 12'hFB2;
iconPixArray[687] = 12'hB81;
iconPixArray[688] = 12'hDA1;
iconPixArray[689] = 12'hFC2;
iconPixArray[690] = 12'hF71;
iconPixArray[691] = 12'h400;
iconPixArray[692] = 12'h567;
iconPixArray[693] = 12'h766;
iconPixArray[694] = 12'h 00;
iconPixArray[695] = 12'h 00;
iconPixArray[696] = 12'h 00;
iconPixArray[697] = 12'h 00;
iconPixArray[698] = 12'h 00;
iconPixArray[699] = 12'h 00;
iconPixArray[700] = 12'h 00;
iconPixArray[701] = 12'h 00;
iconPixArray[702] = 12'h 00;
iconPixArray[703] = 12'h 00;
iconPixArray[704] = 12'h 00;
iconPixArray[705] = 12'h 00;
iconPixArray[706] = 12'h 00;
iconPixArray[707] = 12'h 00;
iconPixArray[708] = 12'h 00;
iconPixArray[709] = 12'h 00;
iconPixArray[710] = 12'h 00;
iconPixArray[711] = 12'h 00;
iconPixArray[712] = 12'h 00;
iconPixArray[713] = 12'h 00;
iconPixArray[714] = 12'h 00;
iconPixArray[715] = 12'h500;
iconPixArray[716] = 12'hF70;
iconPixArray[717] = 12'hE70;
iconPixArray[718] = 12'hF81;
iconPixArray[719] = 12'hFC2;
iconPixArray[720] = 12'hFB2;
iconPixArray[721] = 12'hEC2;
iconPixArray[722] = 12'hE91;
iconPixArray[723] = 12'h710;
iconPixArray[724] = 12'h 00;
iconPixArray[725] = 12'h100;
iconPixArray[726] = 12'h 00;
iconPixArray[727] = 12'h 00;
iconPixArray[728] = 12'h 00;
iconPixArray[729] = 12'h 00;
iconPixArray[730] = 12'h 00;
iconPixArray[731] = 12'h 00;
iconPixArray[732] = 12'h 00;
iconPixArray[733] = 12'h 00;
iconPixArray[734] = 12'h 00;
iconPixArray[735] = 12'h 00;
iconPixArray[736] = 12'h 00;
iconPixArray[737] = 12'h 00;
iconPixArray[738] = 12'h 00;
iconPixArray[739] = 12'h 00;
iconPixArray[740] = 12'h 00;
iconPixArray[741] = 12'h 00;
iconPixArray[742] = 12'h 00;
iconPixArray[743] = 12'h 00;
iconPixArray[744] = 12'h 00;
iconPixArray[745] = 12'h 00;
iconPixArray[746] = 12'h 00;
iconPixArray[747] = 12'hB30;
iconPixArray[748] = 12'hE40;
iconPixArray[749] = 12'hE20;
iconPixArray[750] = 12'hF81;
iconPixArray[751] = 12'hE81;
iconPixArray[752] = 12'hEA1;
iconPixArray[753] = 12'hE60;
iconPixArray[754] = 12'hE71;
iconPixArray[755] = 12'hA20;
iconPixArray[756] = 12'h 00;
iconPixArray[757] = 12'h 00;
iconPixArray[758] = 12'h 00;
iconPixArray[759] = 12'h 00;
iconPixArray[760] = 12'h 00;
iconPixArray[761] = 12'h 00;
iconPixArray[762] = 12'h 00;
iconPixArray[763] = 12'h 00;
iconPixArray[764] = 12'h 00;
iconPixArray[765] = 12'h 00;
iconPixArray[766] = 12'h 00;
iconPixArray[767] = 12'h 00;
iconPixArray[768] = 12'h 00;
iconPixArray[769] = 12'h 00;
iconPixArray[770] = 12'h 00;
iconPixArray[771] = 12'h 00;
iconPixArray[772] = 12'h 00;
iconPixArray[773] = 12'h 00;
iconPixArray[774] = 12'h 00;
iconPixArray[775] = 12'h 00;
iconPixArray[776] = 12'h 00;
iconPixArray[777] = 12'h 00;
iconPixArray[778] = 12'h100;
iconPixArray[779] = 12'hE30;
iconPixArray[780] = 12'hF30;
iconPixArray[781] = 12'hE30;
iconPixArray[782] = 12'hF60;
iconPixArray[783] = 12'hE50;
iconPixArray[784] = 12'hF60;
iconPixArray[785] = 12'hE30;
iconPixArray[786] = 12'hF30;
iconPixArray[787] = 12'hB20;
iconPixArray[788] = 12'h 00;
iconPixArray[789] = 12'h 00;
iconPixArray[790] = 12'h 00;
iconPixArray[791] = 12'h 00;
iconPixArray[792] = 12'h 00;
iconPixArray[793] = 12'h 00;
iconPixArray[794] = 12'h 00;
iconPixArray[795] = 12'h 00;
iconPixArray[796] = 12'h 00;
iconPixArray[797] = 12'h 00;
iconPixArray[798] = 12'h 00;
iconPixArray[799] = 12'h 00;
iconPixArray[800] = 12'h 00;
iconPixArray[801] = 12'h 00;
iconPixArray[802] = 12'h 00;
iconPixArray[803] = 12'h 00;
iconPixArray[804] = 12'h 00;
iconPixArray[805] = 12'h 00;
iconPixArray[806] = 12'h 00;
iconPixArray[807] = 12'h 00;
iconPixArray[808] = 12'h 00;
iconPixArray[809] = 12'h 00;
iconPixArray[810] = 12'h100;
iconPixArray[811] = 12'hB20;
iconPixArray[812] = 12'h820;
iconPixArray[813] = 12'hF30;
iconPixArray[814] = 12'hF30;
iconPixArray[815] = 12'hF30;
iconPixArray[816] = 12'hF30;
iconPixArray[817] = 12'h820;
iconPixArray[818] = 12'hC30;
iconPixArray[819] = 12'hD30;
iconPixArray[820] = 12'h 00;
iconPixArray[821] = 12'h 00;
iconPixArray[822] = 12'h 00;
iconPixArray[823] = 12'h 00;
iconPixArray[824] = 12'h 00;
iconPixArray[825] = 12'h 00;
iconPixArray[826] = 12'h 00;
iconPixArray[827] = 12'h 00;
iconPixArray[828] = 12'h 00;
iconPixArray[829] = 12'h 00;
iconPixArray[830] = 12'h 00;
iconPixArray[831] = 12'h 00;
iconPixArray[832] = 12'h 00;
iconPixArray[833] = 12'h 00;
iconPixArray[834] = 12'h 00;
iconPixArray[835] = 12'h 00;
iconPixArray[836] = 12'h 00;
iconPixArray[837] = 12'h 00;
iconPixArray[838] = 12'h 00;
iconPixArray[839] = 12'h 00;
iconPixArray[840] = 12'h 00;
iconPixArray[841] = 12'h 00;
iconPixArray[842] = 12'h 00;
iconPixArray[843] = 12'h 00;
iconPixArray[844] = 12'h410;
iconPixArray[845] = 12'hE40;
iconPixArray[846] = 12'hD30;
iconPixArray[847] = 12'h920;
iconPixArray[848] = 12'hF40;
iconPixArray[849] = 12'h510;
iconPixArray[850] = 12'h200;
iconPixArray[851] = 12'h820;
iconPixArray[852] = 12'h 00;
iconPixArray[853] = 12'h 00;
iconPixArray[854] = 12'h 00;
iconPixArray[855] = 12'h 00;
iconPixArray[856] = 12'h 00;
iconPixArray[857] = 12'h 00;
iconPixArray[858] = 12'h 00;
iconPixArray[859] = 12'h 00;
iconPixArray[860] = 12'h 00;
iconPixArray[861] = 12'h 00;
iconPixArray[862] = 12'h 00;
iconPixArray[863] = 12'h 00;
iconPixArray[864] = 12'h 00;
iconPixArray[865] = 12'h 00;
iconPixArray[866] = 12'h 00;
iconPixArray[867] = 12'h 00;
iconPixArray[868] = 12'h 00;
iconPixArray[869] = 12'h 00;
iconPixArray[870] = 12'h 00;
iconPixArray[871] = 12'h 00;
iconPixArray[872] = 12'h 00;
iconPixArray[873] = 12'h 00;
iconPixArray[874] = 12'h 00;
iconPixArray[875] = 12'h 00;
iconPixArray[876] = 12'h300;
iconPixArray[877] = 12'hF40;
iconPixArray[878] = 12'h920;
iconPixArray[879] = 12'h 00;
iconPixArray[880] = 12'hE30;
iconPixArray[881] = 12'h610;
iconPixArray[882] = 12'h 00;
iconPixArray[883] = 12'h 00;
iconPixArray[884] = 12'h 00;
iconPixArray[885] = 12'h 00;
iconPixArray[886] = 12'h 00;
iconPixArray[887] = 12'h 00;
iconPixArray[888] = 12'h 00;
iconPixArray[889] = 12'h 00;
iconPixArray[890] = 12'h 00;
iconPixArray[891] = 12'h 00;
iconPixArray[892] = 12'h 00;
iconPixArray[893] = 12'h 00;
iconPixArray[894] = 12'h 00;
iconPixArray[895] = 12'h 00;
iconPixArray[896] = 12'h 00;
iconPixArray[897] = 12'h 00;
iconPixArray[898] = 12'h 00;
iconPixArray[899] = 12'h 00;
iconPixArray[900] = 12'h 00;
iconPixArray[901] = 12'h 00;
iconPixArray[902] = 12'h 00;
iconPixArray[903] = 12'h 00;
iconPixArray[904] = 12'h 00;
iconPixArray[905] = 12'h 00;
iconPixArray[906] = 12'h 00;
iconPixArray[907] = 12'h 00;
iconPixArray[908] = 12'h100;
iconPixArray[909] = 12'hE30;
iconPixArray[910] = 12'h300;
iconPixArray[911] = 12'h 00;
iconPixArray[912] = 12'h820;
iconPixArray[913] = 12'h510;
iconPixArray[914] = 12'h 00;
iconPixArray[915] = 12'h 00;
iconPixArray[916] = 12'h 00;
iconPixArray[917] = 12'h 00;
iconPixArray[918] = 12'h 00;
iconPixArray[919] = 12'h 00;
iconPixArray[920] = 12'h 00;
iconPixArray[921] = 12'h 00;
iconPixArray[922] = 12'h 00;
iconPixArray[923] = 12'h 00;
iconPixArray[924] = 12'h 00;
iconPixArray[925] = 12'h 00;
iconPixArray[926] = 12'h 00;
iconPixArray[927] = 12'h 00;
iconPixArray[928] = 12'h 00;
iconPixArray[929] = 12'h 00;
iconPixArray[930] = 12'h 00;
iconPixArray[931] = 12'h 00;
iconPixArray[932] = 12'h 00;
iconPixArray[933] = 12'h 00;
iconPixArray[934] = 12'h 00;
iconPixArray[935] = 12'h 00;
iconPixArray[936] = 12'h 00;
iconPixArray[937] = 12'h 00;
iconPixArray[938] = 12'h 00;
iconPixArray[939] = 12'h 00;
iconPixArray[940] = 12'h 00;
iconPixArray[941] = 12'h200;
iconPixArray[942] = 12'h 00;
iconPixArray[943] = 12'h 00;
iconPixArray[944] = 12'h 00;
iconPixArray[945] = 12'h 00;
iconPixArray[946] = 12'h 00;
iconPixArray[947] = 12'h 00;
iconPixArray[948] = 12'h 00;
iconPixArray[949] = 12'h 00;
iconPixArray[950] = 12'h 00;
iconPixArray[951] = 12'h 00;
iconPixArray[952] = 12'h 00;
iconPixArray[953] = 12'h 00;
iconPixArray[954] = 12'h 00;
iconPixArray[955] = 12'h 00;
iconPixArray[956] = 12'h 00;
iconPixArray[957] = 12'h 00;
iconPixArray[958] = 12'h 00;
iconPixArray[959] = 12'h 00;
iconPixArray[960] = 12'h 00;
iconPixArray[961] = 12'h 00;
iconPixArray[962] = 12'h 00;
iconPixArray[963] = 12'h 00;
iconPixArray[964] = 12'h 00;
iconPixArray[965] = 12'h 00;
iconPixArray[966] = 12'h 00;
iconPixArray[967] = 12'h 00;
iconPixArray[968] = 12'h 00;
iconPixArray[969] = 12'h 00;
iconPixArray[970] = 12'h 00;
iconPixArray[971] = 12'h 00;
iconPixArray[972] = 12'h 00;
iconPixArray[973] = 12'h 00;
iconPixArray[974] = 12'h 00;
iconPixArray[975] = 12'h 00;
iconPixArray[976] = 12'h 00;
iconPixArray[977] = 12'h 00;
iconPixArray[978] = 12'h 00;
iconPixArray[979] = 12'h 00;
iconPixArray[980] = 12'h 00;
iconPixArray[981] = 12'h 00;
iconPixArray[982] = 12'h 00;
iconPixArray[983] = 12'h 00;
iconPixArray[984] = 12'h 00;
iconPixArray[985] = 12'h 00;
iconPixArray[986] = 12'h 00;
iconPixArray[987] = 12'h 00;
iconPixArray[988] = 12'h 00;
iconPixArray[989] = 12'h 00;
iconPixArray[990] = 12'h 00;
iconPixArray[991] = 12'h 00;
iconPixArray[992] = 12'h 00;
iconPixArray[993] = 12'h 00;
iconPixArray[994] = 12'h 00;
iconPixArray[995] = 12'h 00;
iconPixArray[996] = 12'h 00;
iconPixArray[997] = 12'h 00;
iconPixArray[998] = 12'h 00;
iconPixArray[999] = 12'h 00;
iconPixArray[1000] = 12'h 00;
iconPixArray[1001] = 12'h 00;
iconPixArray[1002] = 12'h 00;
iconPixArray[1003] = 12'h 00;
iconPixArray[1004] = 12'h 00;
iconPixArray[1005] = 12'h 00;
iconPixArray[1006] = 12'h 00;
iconPixArray[1007] = 12'h 00;
iconPixArray[1008] = 12'h 00;
iconPixArray[1009] = 12'h 00;
iconPixArray[1010] = 12'h 00;
iconPixArray[1011] = 12'h 00;
iconPixArray[1012] = 12'h 00;
iconPixArray[1013] = 12'h 00;
iconPixArray[1014] = 12'h 00;
iconPixArray[1015] = 12'h 00;
iconPixArray[1016] = 12'h 00;
iconPixArray[1017] = 12'h 00;
iconPixArray[1018] = 12'h 00;
iconPixArray[1019] = 12'h 00;
iconPixArray[1020] = 12'h 00;
iconPixArray[1021] = 12'h 00;
iconPixArray[1022] = 12'h 00;
iconPixArray[1023] = 12'h 00;
iconPixArray[1024] = 12'h 00;
iconPixArray[1025] = 12'h 00;
iconPixArray[1026] = 12'h 00;
iconPixArray[1027] = 12'h 00;
iconPixArray[1028] = 12'h 00;
iconPixArray[1029] = 12'h 00;
iconPixArray[1030] = 12'h 00;
iconPixArray[1031] = 12'h 00;
iconPixArray[1032] = 12'h 00;
iconPixArray[1033] = 12'h 00;
iconPixArray[1034] = 12'h 00;
iconPixArray[1035] = 12'h 00;
iconPixArray[1036] = 12'h 00;
iconPixArray[1037] = 12'h 00;
iconPixArray[1038] = 12'h 00;
iconPixArray[1039] = 12'h 00;
iconPixArray[1040] = 12'h 00;
iconPixArray[1041] = 12'h 00;
iconPixArray[1042] = 12'h 00;
iconPixArray[1043] = 12'h 00;
iconPixArray[1044] = 12'h 00;
iconPixArray[1045] = 12'h 00;
iconPixArray[1046] = 12'h 00;
iconPixArray[1047] = 12'h 00;
iconPixArray[1048] = 12'h 00;
iconPixArray[1049] = 12'h 00;
iconPixArray[1050] = 12'h 00;
iconPixArray[1051] = 12'h 00;
iconPixArray[1052] = 12'h 00;
iconPixArray[1053] = 12'h 00;
iconPixArray[1054] = 12'h 00;
iconPixArray[1055] = 12'h 00;
iconPixArray[1056] = 12'h 00;
iconPixArray[1057] = 12'h 00;
iconPixArray[1058] = 12'h 00;
iconPixArray[1059] = 12'h 00;
iconPixArray[1060] = 12'h 00;
iconPixArray[1061] = 12'h 00;
iconPixArray[1062] = 12'h 00;
iconPixArray[1063] = 12'h 00;
iconPixArray[1064] = 12'h 00;
iconPixArray[1065] = 12'h 00;
iconPixArray[1066] = 12'h 00;
iconPixArray[1067] = 12'h 00;
iconPixArray[1068] = 12'h 00;
iconPixArray[1069] = 12'h 00;
iconPixArray[1070] = 12'h 00;
iconPixArray[1071] = 12'h 00;
iconPixArray[1072] = 12'h 00;
iconPixArray[1073] = 12'h 00;
iconPixArray[1074] = 12'h 00;
iconPixArray[1075] = 12'h 00;
iconPixArray[1076] = 12'h 00;
iconPixArray[1077] = 12'h 00;
iconPixArray[1078] = 12'h 00;
iconPixArray[1079] = 12'h 00;
iconPixArray[1080] = 12'h 00;
iconPixArray[1081] = 12'h 00;
iconPixArray[1082] = 12'h 00;
iconPixArray[1083] = 12'h 00;
iconPixArray[1084] = 12'h 00;
iconPixArray[1085] = 12'h 00;
iconPixArray[1086] = 12'h 00;
iconPixArray[1087] = 12'h 00;
iconPixArray[1088] = 12'h 00;
iconPixArray[1089] = 12'h 00;
iconPixArray[1090] = 12'h 00;
iconPixArray[1091] = 12'h 00;
iconPixArray[1092] = 12'h 00;
iconPixArray[1093] = 12'h 00;
iconPixArray[1094] = 12'h 00;
iconPixArray[1095] = 12'h 00;
iconPixArray[1096] = 12'h 00;
iconPixArray[1097] = 12'h 00;
iconPixArray[1098] = 12'h 00;
iconPixArray[1099] = 12'h 00;
iconPixArray[1100] = 12'h 00;
iconPixArray[1101] = 12'h 00;
iconPixArray[1102] = 12'h 00;
iconPixArray[1103] = 12'h333;
iconPixArray[1104] = 12'h999;
iconPixArray[1105] = 12'h 00;
iconPixArray[1106] = 12'h 00;
iconPixArray[1107] = 12'h 00;
iconPixArray[1108] = 12'h 00;
iconPixArray[1109] = 12'h 00;
iconPixArray[1110] = 12'h 00;
iconPixArray[1111] = 12'h 00;
iconPixArray[1112] = 12'h 00;
iconPixArray[1113] = 12'h 00;
iconPixArray[1114] = 12'h 00;
iconPixArray[1115] = 12'h 00;
iconPixArray[1116] = 12'h 00;
iconPixArray[1117] = 12'h 00;
iconPixArray[1118] = 12'h 00;
iconPixArray[1119] = 12'h 00;
iconPixArray[1120] = 12'h 00;
iconPixArray[1121] = 12'h 00;
iconPixArray[1122] = 12'h 00;
iconPixArray[1123] = 12'h 00;
iconPixArray[1124] = 12'h 00;
iconPixArray[1125] = 12'h 00;
iconPixArray[1126] = 12'h 00;
iconPixArray[1127] = 12'h 00;
iconPixArray[1128] = 12'h 00;
iconPixArray[1129] = 12'h 00;
iconPixArray[1130] = 12'h 00;
iconPixArray[1131] = 12'h 00;
iconPixArray[1132] = 12'h 00;
iconPixArray[1133] = 12'h 00;
iconPixArray[1134] = 12'h 00;
iconPixArray[1135] = 12'hBBB;
iconPixArray[1136] = 12'hEEE;
iconPixArray[1137] = 12'h666;
iconPixArray[1138] = 12'h 00;
iconPixArray[1139] = 12'h 00;
iconPixArray[1140] = 12'h 00;
iconPixArray[1141] = 12'h 00;
iconPixArray[1142] = 12'h 00;
iconPixArray[1143] = 12'h 00;
iconPixArray[1144] = 12'h 00;
iconPixArray[1145] = 12'h 00;
iconPixArray[1146] = 12'h 00;
iconPixArray[1147] = 12'h 00;
iconPixArray[1148] = 12'h 00;
iconPixArray[1149] = 12'h 00;
iconPixArray[1150] = 12'h 00;
iconPixArray[1151] = 12'h 00;
iconPixArray[1152] = 12'h 00;
iconPixArray[1153] = 12'h 00;
iconPixArray[1154] = 12'h 00;
iconPixArray[1155] = 12'h 00;
iconPixArray[1156] = 12'h 00;
iconPixArray[1157] = 12'h 00;
iconPixArray[1158] = 12'h 00;
iconPixArray[1159] = 12'h 00;
iconPixArray[1160] = 12'h 00;
iconPixArray[1161] = 12'h 00;
iconPixArray[1162] = 12'h 00;
iconPixArray[1163] = 12'h 00;
iconPixArray[1164] = 12'h 00;
iconPixArray[1165] = 12'h 00;
iconPixArray[1166] = 12'h666;
iconPixArray[1167] = 12'hDDD;
iconPixArray[1168] = 12'hCCC;
iconPixArray[1169] = 12'hCCC;
iconPixArray[1170] = 12'h222;
iconPixArray[1171] = 12'h 00;
iconPixArray[1172] = 12'h 00;
iconPixArray[1173] = 12'h 00;
iconPixArray[1174] = 12'h 00;
iconPixArray[1175] = 12'h 00;
iconPixArray[1176] = 12'h 00;
iconPixArray[1177] = 12'h 00;
iconPixArray[1178] = 12'h 00;
iconPixArray[1179] = 12'h 00;
iconPixArray[1180] = 12'h 00;
iconPixArray[1181] = 12'h 00;
iconPixArray[1182] = 12'h 00;
iconPixArray[1183] = 12'h 00;
iconPixArray[1184] = 12'h 00;
iconPixArray[1185] = 12'h 00;
iconPixArray[1186] = 12'h 00;
iconPixArray[1187] = 12'h 00;
iconPixArray[1188] = 12'h 00;
iconPixArray[1189] = 12'h 00;
iconPixArray[1190] = 12'h 00;
iconPixArray[1191] = 12'h 00;
iconPixArray[1192] = 12'h 00;
iconPixArray[1193] = 12'h 00;
iconPixArray[1194] = 12'h 00;
iconPixArray[1195] = 12'h 00;
iconPixArray[1196] = 12'h 00;
iconPixArray[1197] = 12'h111;
iconPixArray[1198] = 12'hCCC;
iconPixArray[1199] = 12'hCCC;
iconPixArray[1200] = 12'hCCC;
iconPixArray[1201] = 12'hDDD;
iconPixArray[1202] = 12'h888;
iconPixArray[1203] = 12'h 00;
iconPixArray[1204] = 12'h 00;
iconPixArray[1205] = 12'h 00;
iconPixArray[1206] = 12'h 00;
iconPixArray[1207] = 12'h 00;
iconPixArray[1208] = 12'h 00;
iconPixArray[1209] = 12'h 00;
iconPixArray[1210] = 12'h 00;
iconPixArray[1211] = 12'h 00;
iconPixArray[1212] = 12'h 00;
iconPixArray[1213] = 12'h 00;
iconPixArray[1214] = 12'h 00;
iconPixArray[1215] = 12'h 00;
iconPixArray[1216] = 12'h 00;
iconPixArray[1217] = 12'h 00;
iconPixArray[1218] = 12'h 00;
iconPixArray[1219] = 12'h 00;
iconPixArray[1220] = 12'h 00;
iconPixArray[1221] = 12'h 00;
iconPixArray[1222] = 12'h 00;
iconPixArray[1223] = 12'h 00;
iconPixArray[1224] = 12'h 00;
iconPixArray[1225] = 12'h 00;
iconPixArray[1226] = 12'h 00;
iconPixArray[1227] = 12'h 00;
iconPixArray[1228] = 12'h 00;
iconPixArray[1229] = 12'h666;
iconPixArray[1230] = 12'hDDD;
iconPixArray[1231] = 12'hCCC;
iconPixArray[1232] = 12'hDDD;
iconPixArray[1233] = 12'hCCC;
iconPixArray[1234] = 12'hDDD;
iconPixArray[1235] = 12'h222;
iconPixArray[1236] = 12'h 00;
iconPixArray[1237] = 12'h 00;
iconPixArray[1238] = 12'h 00;
iconPixArray[1239] = 12'h 00;
iconPixArray[1240] = 12'h 00;
iconPixArray[1241] = 12'h 00;
iconPixArray[1242] = 12'h 00;
iconPixArray[1243] = 12'h 00;
iconPixArray[1244] = 12'h 00;
iconPixArray[1245] = 12'h 00;
iconPixArray[1246] = 12'h 00;
iconPixArray[1247] = 12'h 00;
iconPixArray[1248] = 12'h 00;
iconPixArray[1249] = 12'h 00;
iconPixArray[1250] = 12'h 00;
iconPixArray[1251] = 12'h 00;
iconPixArray[1252] = 12'h 00;
iconPixArray[1253] = 12'h 00;
iconPixArray[1254] = 12'h 00;
iconPixArray[1255] = 12'h 00;
iconPixArray[1256] = 12'h 00;
iconPixArray[1257] = 12'h 00;
iconPixArray[1258] = 12'h 00;
iconPixArray[1259] = 12'h 00;
iconPixArray[1260] = 12'h 00;
iconPixArray[1261] = 12'hAAA;
iconPixArray[1262] = 12'hDDD;
iconPixArray[1263] = 12'hCCC;
iconPixArray[1264] = 12'hBBB;
iconPixArray[1265] = 12'hDDD;
iconPixArray[1266] = 12'hDDD;
iconPixArray[1267] = 12'h777;
iconPixArray[1268] = 12'h 00;
iconPixArray[1269] = 12'h 00;
iconPixArray[1270] = 12'h 00;
iconPixArray[1271] = 12'h 00;
iconPixArray[1272] = 12'h 00;
iconPixArray[1273] = 12'h 00;
iconPixArray[1274] = 12'h 00;
iconPixArray[1275] = 12'h 00;
iconPixArray[1276] = 12'h 00;
iconPixArray[1277] = 12'h 00;
iconPixArray[1278] = 12'h 00;
iconPixArray[1279] = 12'h 00;
iconPixArray[1280] = 12'h 00;
iconPixArray[1281] = 12'h 00;
iconPixArray[1282] = 12'h 00;
iconPixArray[1283] = 12'h 00;
iconPixArray[1284] = 12'h 00;
iconPixArray[1285] = 12'h 00;
iconPixArray[1286] = 12'h 00;
iconPixArray[1287] = 12'h 00;
iconPixArray[1288] = 12'h 00;
iconPixArray[1289] = 12'h 00;
iconPixArray[1290] = 12'h 00;
iconPixArray[1291] = 12'h 00;
iconPixArray[1292] = 12'h222;
iconPixArray[1293] = 12'hDDD;
iconPixArray[1294] = 12'hAAA;
iconPixArray[1295] = 12'h222;
iconPixArray[1296] = 12'h222;
iconPixArray[1297] = 12'h666;
iconPixArray[1298] = 12'hDDD;
iconPixArray[1299] = 12'hBBB;
iconPixArray[1300] = 12'h 00;
iconPixArray[1301] = 12'h 00;
iconPixArray[1302] = 12'h 00;
iconPixArray[1303] = 12'h 00;
iconPixArray[1304] = 12'h 00;
iconPixArray[1305] = 12'h 00;
iconPixArray[1306] = 12'h 00;
iconPixArray[1307] = 12'h 00;
iconPixArray[1308] = 12'h 00;
iconPixArray[1309] = 12'h 00;
iconPixArray[1310] = 12'h 00;
iconPixArray[1311] = 12'h 00;
iconPixArray[1312] = 12'h 00;
iconPixArray[1313] = 12'h 00;
iconPixArray[1314] = 12'h 00;
iconPixArray[1315] = 12'h 00;
iconPixArray[1316] = 12'h 00;
iconPixArray[1317] = 12'h 00;
iconPixArray[1318] = 12'h 00;
iconPixArray[1319] = 12'h 00;
iconPixArray[1320] = 12'h 00;
iconPixArray[1321] = 12'h 00;
iconPixArray[1322] = 12'h 00;
iconPixArray[1323] = 12'h 00;
iconPixArray[1324] = 12'h444;
iconPixArray[1325] = 12'hEEE;
iconPixArray[1326] = 12'h444;
iconPixArray[1327] = 12'h799;
iconPixArray[1328] = 12'hBDD;
iconPixArray[1329] = 12'h222;
iconPixArray[1330] = 12'hAAA;
iconPixArray[1331] = 12'hDDD;
iconPixArray[1332] = 12'h333;
iconPixArray[1333] = 12'h 00;
iconPixArray[1334] = 12'h 00;
iconPixArray[1335] = 12'h 00;
iconPixArray[1336] = 12'h 00;
iconPixArray[1337] = 12'h 00;
iconPixArray[1338] = 12'h 00;
iconPixArray[1339] = 12'h 00;
iconPixArray[1340] = 12'h 00;
iconPixArray[1341] = 12'h 00;
iconPixArray[1342] = 12'h 00;
iconPixArray[1343] = 12'h 00;
iconPixArray[1344] = 12'h 00;
iconPixArray[1345] = 12'h 00;
iconPixArray[1346] = 12'h 00;
iconPixArray[1347] = 12'h 00;
iconPixArray[1348] = 12'h 00;
iconPixArray[1349] = 12'h 00;
iconPixArray[1350] = 12'h 00;
iconPixArray[1351] = 12'h 00;
iconPixArray[1352] = 12'h 00;
iconPixArray[1353] = 12'h 00;
iconPixArray[1354] = 12'h 00;
iconPixArray[1355] = 12'h 00;
iconPixArray[1356] = 12'h777;
iconPixArray[1357] = 12'hEEE;
iconPixArray[1358] = 12'h444;
iconPixArray[1359] = 12'h688;
iconPixArray[1360] = 12'hBDD;
iconPixArray[1361] = 12'h222;
iconPixArray[1362] = 12'hAAA;
iconPixArray[1363] = 12'hEEE;
iconPixArray[1364] = 12'h666;
iconPixArray[1365] = 12'h 00;
iconPixArray[1366] = 12'h 00;
iconPixArray[1367] = 12'h 00;
iconPixArray[1368] = 12'h 00;
iconPixArray[1369] = 12'h 00;
iconPixArray[1370] = 12'h 00;
iconPixArray[1371] = 12'h 00;
iconPixArray[1372] = 12'h 00;
iconPixArray[1373] = 12'h 00;
iconPixArray[1374] = 12'h 00;
iconPixArray[1375] = 12'h 00;
iconPixArray[1376] = 12'h 00;
iconPixArray[1377] = 12'h 00;
iconPixArray[1378] = 12'h 00;
iconPixArray[1379] = 12'h 00;
iconPixArray[1380] = 12'h 00;
iconPixArray[1381] = 12'h 00;
iconPixArray[1382] = 12'h 00;
iconPixArray[1383] = 12'h 00;
iconPixArray[1384] = 12'h 00;
iconPixArray[1385] = 12'h 00;
iconPixArray[1386] = 12'h 00;
iconPixArray[1387] = 12'h 00;
iconPixArray[1388] = 12'h888;
iconPixArray[1389] = 12'hEEE;
iconPixArray[1390] = 12'hAAA;
iconPixArray[1391] = 12'h222;
iconPixArray[1392] = 12'h222;
iconPixArray[1393] = 12'h666;
iconPixArray[1394] = 12'hDDD;
iconPixArray[1395] = 12'hDDD;
iconPixArray[1396] = 12'h888;
iconPixArray[1397] = 12'h 00;
iconPixArray[1398] = 12'h 00;
iconPixArray[1399] = 12'h 00;
iconPixArray[1400] = 12'h 00;
iconPixArray[1401] = 12'h 00;
iconPixArray[1402] = 12'h 00;
iconPixArray[1403] = 12'h 00;
iconPixArray[1404] = 12'h 00;
iconPixArray[1405] = 12'h 00;
iconPixArray[1406] = 12'h 00;
iconPixArray[1407] = 12'h 00;
iconPixArray[1408] = 12'h 00;
iconPixArray[1409] = 12'h 00;
iconPixArray[1410] = 12'h 00;
iconPixArray[1411] = 12'h 00;
iconPixArray[1412] = 12'h 00;
iconPixArray[1413] = 12'h 00;
iconPixArray[1414] = 12'h 00;
iconPixArray[1415] = 12'h 00;
iconPixArray[1416] = 12'h 00;
iconPixArray[1417] = 12'h 00;
iconPixArray[1418] = 12'h 00;
iconPixArray[1419] = 12'h 00;
iconPixArray[1420] = 12'h999;
iconPixArray[1421] = 12'hDDD;
iconPixArray[1422] = 12'hDDD;
iconPixArray[1423] = 12'hCCC;
iconPixArray[1424] = 12'hBBB;
iconPixArray[1425] = 12'hDDD;
iconPixArray[1426] = 12'hCCC;
iconPixArray[1427] = 12'hDDD;
iconPixArray[1428] = 12'h999;
iconPixArray[1429] = 12'h 00;
iconPixArray[1430] = 12'h 00;
iconPixArray[1431] = 12'h 00;
iconPixArray[1432] = 12'h 00;
iconPixArray[1433] = 12'h 00;
iconPixArray[1434] = 12'h 00;
iconPixArray[1435] = 12'h 00;
iconPixArray[1436] = 12'h 00;
iconPixArray[1437] = 12'h 00;
iconPixArray[1438] = 12'h 00;
iconPixArray[1439] = 12'h 00;
iconPixArray[1440] = 12'h 00;
iconPixArray[1441] = 12'h 00;
iconPixArray[1442] = 12'h 00;
iconPixArray[1443] = 12'h 00;
iconPixArray[1444] = 12'h 00;
iconPixArray[1445] = 12'h 00;
iconPixArray[1446] = 12'h 00;
iconPixArray[1447] = 12'h 00;
iconPixArray[1448] = 12'h 00;
iconPixArray[1449] = 12'h 00;
iconPixArray[1450] = 12'h 00;
iconPixArray[1451] = 12'h 00;
iconPixArray[1452] = 12'hAAA;
iconPixArray[1453] = 12'hDDD;
iconPixArray[1454] = 12'hCCC;
iconPixArray[1455] = 12'hCCC;
iconPixArray[1456] = 12'hCCC;
iconPixArray[1457] = 12'hCCC;
iconPixArray[1458] = 12'hCCC;
iconPixArray[1459] = 12'hDDD;
iconPixArray[1460] = 12'h999;
iconPixArray[1461] = 12'h 00;
iconPixArray[1462] = 12'h 00;
iconPixArray[1463] = 12'h 00;
iconPixArray[1464] = 12'h 00;
iconPixArray[1465] = 12'h 00;
iconPixArray[1466] = 12'h 00;
iconPixArray[1467] = 12'h 00;
iconPixArray[1468] = 12'h 00;
iconPixArray[1469] = 12'h 00;
iconPixArray[1470] = 12'h 00;
iconPixArray[1471] = 12'h 00;
iconPixArray[1472] = 12'h 00;
iconPixArray[1473] = 12'h 00;
iconPixArray[1474] = 12'h 00;
iconPixArray[1475] = 12'h 00;
iconPixArray[1476] = 12'h 00;
iconPixArray[1477] = 12'h 00;
iconPixArray[1478] = 12'h 00;
iconPixArray[1479] = 12'h 00;
iconPixArray[1480] = 12'h 00;
iconPixArray[1481] = 12'h 00;
iconPixArray[1482] = 12'h 00;
iconPixArray[1483] = 12'h 00;
iconPixArray[1484] = 12'hAAA;
iconPixArray[1485] = 12'hDDD;
iconPixArray[1486] = 12'hCCC;
iconPixArray[1487] = 12'h666;
iconPixArray[1488] = 12'h333;
iconPixArray[1489] = 12'hAAA;
iconPixArray[1490] = 12'hDDD;
iconPixArray[1491] = 12'hDDD;
iconPixArray[1492] = 12'h999;
iconPixArray[1493] = 12'h 00;
iconPixArray[1494] = 12'h 00;
iconPixArray[1495] = 12'h 00;
iconPixArray[1496] = 12'h 00;
iconPixArray[1497] = 12'h 00;
iconPixArray[1498] = 12'h 00;
iconPixArray[1499] = 12'h 00;
iconPixArray[1500] = 12'h 00;
iconPixArray[1501] = 12'h 00;
iconPixArray[1502] = 12'h 00;
iconPixArray[1503] = 12'h 00;
iconPixArray[1504] = 12'h 00;
iconPixArray[1505] = 12'h 00;
iconPixArray[1506] = 12'h 00;
iconPixArray[1507] = 12'h 00;
iconPixArray[1508] = 12'h 00;
iconPixArray[1509] = 12'h 00;
iconPixArray[1510] = 12'h 00;
iconPixArray[1511] = 12'h 00;
iconPixArray[1512] = 12'h 00;
iconPixArray[1513] = 12'h 00;
iconPixArray[1514] = 12'h111;
iconPixArray[1515] = 12'h555;
iconPixArray[1516] = 12'h999;
iconPixArray[1517] = 12'hEEE;
iconPixArray[1518] = 12'hAAA;
iconPixArray[1519] = 12'h666;
iconPixArray[1520] = 12'h333;
iconPixArray[1521] = 12'hAAA;
iconPixArray[1522] = 12'hDDD;
iconPixArray[1523] = 12'hDDD;
iconPixArray[1524] = 12'h888;
iconPixArray[1525] = 12'h111;
iconPixArray[1526] = 12'h 00;
iconPixArray[1527] = 12'h 00;
iconPixArray[1528] = 12'h 00;
iconPixArray[1529] = 12'h 00;
iconPixArray[1530] = 12'h 00;
iconPixArray[1531] = 12'h 00;
iconPixArray[1532] = 12'h 00;
iconPixArray[1533] = 12'h 00;
iconPixArray[1534] = 12'h 00;
iconPixArray[1535] = 12'h 00;
iconPixArray[1536] = 12'h 00;
iconPixArray[1537] = 12'h 00;
iconPixArray[1538] = 12'h 00;
iconPixArray[1539] = 12'h 00;
iconPixArray[1540] = 12'h 00;
iconPixArray[1541] = 12'h 00;
iconPixArray[1542] = 12'h 00;
iconPixArray[1543] = 12'h 00;
iconPixArray[1544] = 12'h 00;
iconPixArray[1545] = 12'h111;
iconPixArray[1546] = 12'h999;
iconPixArray[1547] = 12'h999;
iconPixArray[1548] = 12'h888;
iconPixArray[1549] = 12'hEEE;
iconPixArray[1550] = 12'h999;
iconPixArray[1551] = 12'h666;
iconPixArray[1552] = 12'h444;
iconPixArray[1553] = 12'hAAA;
iconPixArray[1554] = 12'hDDD;
iconPixArray[1555] = 12'hDDD;
iconPixArray[1556] = 12'h777;
iconPixArray[1557] = 12'h999;
iconPixArray[1558] = 12'h111;
iconPixArray[1559] = 12'h 00;
iconPixArray[1560] = 12'h 00;
iconPixArray[1561] = 12'h 00;
iconPixArray[1562] = 12'h 00;
iconPixArray[1563] = 12'h 00;
iconPixArray[1564] = 12'h 00;
iconPixArray[1565] = 12'h 00;
iconPixArray[1566] = 12'h 00;
iconPixArray[1567] = 12'h 00;
iconPixArray[1568] = 12'h 00;
iconPixArray[1569] = 12'h 00;
iconPixArray[1570] = 12'h 00;
iconPixArray[1571] = 12'h 00;
iconPixArray[1572] = 12'h 00;
iconPixArray[1573] = 12'h 00;
iconPixArray[1574] = 12'h 00;
iconPixArray[1575] = 12'h 00;
iconPixArray[1576] = 12'h 00;
iconPixArray[1577] = 12'h555;
iconPixArray[1578] = 12'hCCC;
iconPixArray[1579] = 12'h999;
iconPixArray[1580] = 12'h777;
iconPixArray[1581] = 12'hDDD;
iconPixArray[1582] = 12'h999;
iconPixArray[1583] = 12'h666;
iconPixArray[1584] = 12'h444;
iconPixArray[1585] = 12'hAAA;
iconPixArray[1586] = 12'hDDD;
iconPixArray[1587] = 12'hCCC;
iconPixArray[1588] = 12'h666;
iconPixArray[1589] = 12'hBBB;
iconPixArray[1590] = 12'h999;
iconPixArray[1591] = 12'h 00;
iconPixArray[1592] = 12'h 00;
iconPixArray[1593] = 12'h 00;
iconPixArray[1594] = 12'h 00;
iconPixArray[1595] = 12'h 00;
iconPixArray[1596] = 12'h 00;
iconPixArray[1597] = 12'h 00;
iconPixArray[1598] = 12'h 00;
iconPixArray[1599] = 12'h 00;
iconPixArray[1600] = 12'h 00;
iconPixArray[1601] = 12'h 00;
iconPixArray[1602] = 12'h 00;
iconPixArray[1603] = 12'h 00;
iconPixArray[1604] = 12'h 00;
iconPixArray[1605] = 12'h 00;
iconPixArray[1606] = 12'h 00;
iconPixArray[1607] = 12'h 00;
iconPixArray[1608] = 12'h 00;
iconPixArray[1609] = 12'h222;
iconPixArray[1610] = 12'hBBB;
iconPixArray[1611] = 12'hAAA;
iconPixArray[1612] = 12'h666;
iconPixArray[1613] = 12'hEEE;
iconPixArray[1614] = 12'hAAB;
iconPixArray[1615] = 12'h666;
iconPixArray[1616] = 12'h444;
iconPixArray[1617] = 12'hBBB;
iconPixArray[1618] = 12'hEEE;
iconPixArray[1619] = 12'hAAA;
iconPixArray[1620] = 12'h666;
iconPixArray[1621] = 12'hCCC;
iconPixArray[1622] = 12'hAAA;
iconPixArray[1623] = 12'h 00;
iconPixArray[1624] = 12'h 00;
iconPixArray[1625] = 12'h 00;
iconPixArray[1626] = 12'h 00;
iconPixArray[1627] = 12'h 00;
iconPixArray[1628] = 12'h 00;
iconPixArray[1629] = 12'h 00;
iconPixArray[1630] = 12'h 00;
iconPixArray[1631] = 12'h 00;
iconPixArray[1632] = 12'h 00;
iconPixArray[1633] = 12'h 00;
iconPixArray[1634] = 12'h 00;
iconPixArray[1635] = 12'h 00;
iconPixArray[1636] = 12'h 00;
iconPixArray[1637] = 12'h 00;
iconPixArray[1638] = 12'h 00;
iconPixArray[1639] = 12'h 00;
iconPixArray[1640] = 12'h 00;
iconPixArray[1641] = 12'h 00;
iconPixArray[1642] = 12'h999;
iconPixArray[1643] = 12'hCCC;
iconPixArray[1644] = 12'h666;
iconPixArray[1645] = 12'h888;
iconPixArray[1646] = 12'h666;
iconPixArray[1647] = 12'h666;
iconPixArray[1648] = 12'h344;
iconPixArray[1649] = 12'h666;
iconPixArray[1650] = 12'hABB;
iconPixArray[1651] = 12'h677;
iconPixArray[1652] = 12'h999;
iconPixArray[1653] = 12'hCCC;
iconPixArray[1654] = 12'h555;
iconPixArray[1655] = 12'h 00;
iconPixArray[1656] = 12'h 00;
iconPixArray[1657] = 12'h 00;
iconPixArray[1658] = 12'h 00;
iconPixArray[1659] = 12'h 00;
iconPixArray[1660] = 12'h 00;
iconPixArray[1661] = 12'h 00;
iconPixArray[1662] = 12'h 00;
iconPixArray[1663] = 12'h 00;
iconPixArray[1664] = 12'h 00;
iconPixArray[1665] = 12'h 00;
iconPixArray[1666] = 12'h 00;
iconPixArray[1667] = 12'h 00;
iconPixArray[1668] = 12'h 00;
iconPixArray[1669] = 12'h 00;
iconPixArray[1670] = 12'h 00;
iconPixArray[1671] = 12'h 00;
iconPixArray[1672] = 12'h 00;
iconPixArray[1673] = 12'h 00;
iconPixArray[1674] = 12'h777;
iconPixArray[1675] = 12'hBCC;
iconPixArray[1676] = 12'h522;
iconPixArray[1677] = 12'hB50;
iconPixArray[1678] = 12'hB90;
iconPixArray[1679] = 12'h444;
iconPixArray[1680] = 12'h432;
iconPixArray[1681] = 12'hB91;
iconPixArray[1682] = 12'h930;
iconPixArray[1683] = 12'h422;
iconPixArray[1684] = 12'hBBB;
iconPixArray[1685] = 12'hAAA;
iconPixArray[1686] = 12'h111;
iconPixArray[1687] = 12'h 00;
iconPixArray[1688] = 12'h 00;
iconPixArray[1689] = 12'h 00;
iconPixArray[1690] = 12'h 00;
iconPixArray[1691] = 12'h 00;
iconPixArray[1692] = 12'h 00;
iconPixArray[1693] = 12'h 00;
iconPixArray[1694] = 12'h 00;
iconPixArray[1695] = 12'h 00;
iconPixArray[1696] = 12'h 00;
iconPixArray[1697] = 12'h 00;
iconPixArray[1698] = 12'h 00;
iconPixArray[1699] = 12'h 00;
iconPixArray[1700] = 12'h 00;
iconPixArray[1701] = 12'h 00;
iconPixArray[1702] = 12'h 00;
iconPixArray[1703] = 12'h 00;
iconPixArray[1704] = 12'h 00;
iconPixArray[1705] = 12'h 00;
iconPixArray[1706] = 12'h333;
iconPixArray[1707] = 12'h434;
iconPixArray[1708] = 12'hB30;
iconPixArray[1709] = 12'hFC2;
iconPixArray[1710] = 12'hFB2;
iconPixArray[1711] = 12'hB81;
iconPixArray[1712] = 12'hDA1;
iconPixArray[1713] = 12'hFC2;
iconPixArray[1714] = 12'hF71;
iconPixArray[1715] = 12'h400;
iconPixArray[1716] = 12'h567;
iconPixArray[1717] = 12'h766;
iconPixArray[1718] = 12'h 00;
iconPixArray[1719] = 12'h 00;
iconPixArray[1720] = 12'h 00;
iconPixArray[1721] = 12'h 00;
iconPixArray[1722] = 12'h 00;
iconPixArray[1723] = 12'h 00;
iconPixArray[1724] = 12'h 00;
iconPixArray[1725] = 12'h 00;
iconPixArray[1726] = 12'h 00;
iconPixArray[1727] = 12'h 00;
iconPixArray[1728] = 12'h 00;
iconPixArray[1729] = 12'h 00;
iconPixArray[1730] = 12'h 00;
iconPixArray[1731] = 12'h 00;
iconPixArray[1732] = 12'h 00;
iconPixArray[1733] = 12'h 00;
iconPixArray[1734] = 12'h 00;
iconPixArray[1735] = 12'h 00;
iconPixArray[1736] = 12'h 00;
iconPixArray[1737] = 12'h 00;
iconPixArray[1738] = 12'h 00;
iconPixArray[1739] = 12'h500;
iconPixArray[1740] = 12'hF70;
iconPixArray[1741] = 12'hE70;
iconPixArray[1742] = 12'hF81;
iconPixArray[1743] = 12'hFC2;
iconPixArray[1744] = 12'hFB2;
iconPixArray[1745] = 12'hEC2;
iconPixArray[1746] = 12'hE91;
iconPixArray[1747] = 12'h710;
iconPixArray[1748] = 12'h 00;
iconPixArray[1749] = 12'h100;
iconPixArray[1750] = 12'h 00;
iconPixArray[1751] = 12'h 00;
iconPixArray[1752] = 12'h 00;
iconPixArray[1753] = 12'h 00;
iconPixArray[1754] = 12'h 00;
iconPixArray[1755] = 12'h 00;
iconPixArray[1756] = 12'h 00;
iconPixArray[1757] = 12'h 00;
iconPixArray[1758] = 12'h 00;
iconPixArray[1759] = 12'h 00;
iconPixArray[1760] = 12'h 00;
iconPixArray[1761] = 12'h 00;
iconPixArray[1762] = 12'h 00;
iconPixArray[1763] = 12'h 00;
iconPixArray[1764] = 12'h 00;
iconPixArray[1765] = 12'h 00;
iconPixArray[1766] = 12'h 00;
iconPixArray[1767] = 12'h 00;
iconPixArray[1768] = 12'h 00;
iconPixArray[1769] = 12'h 00;
iconPixArray[1770] = 12'h 00;
iconPixArray[1771] = 12'hB30;
iconPixArray[1772] = 12'hE40;
iconPixArray[1773] = 12'hE20;
iconPixArray[1774] = 12'hF81;
iconPixArray[1775] = 12'hE81;
iconPixArray[1776] = 12'hEA1;
iconPixArray[1777] = 12'hE60;
iconPixArray[1778] = 12'hE71;
iconPixArray[1779] = 12'hA20;
iconPixArray[1780] = 12'h 00;
iconPixArray[1781] = 12'h 00;
iconPixArray[1782] = 12'h 00;
iconPixArray[1783] = 12'h 00;
iconPixArray[1784] = 12'h 00;
iconPixArray[1785] = 12'h 00;
iconPixArray[1786] = 12'h 00;
iconPixArray[1787] = 12'h 00;
iconPixArray[1788] = 12'h 00;
iconPixArray[1789] = 12'h 00;
iconPixArray[1790] = 12'h 00;
iconPixArray[1791] = 12'h 00;
iconPixArray[1792] = 12'h 00;
iconPixArray[1793] = 12'h 00;
iconPixArray[1794] = 12'h 00;
iconPixArray[1795] = 12'h 00;
iconPixArray[1796] = 12'h 00;
iconPixArray[1797] = 12'h 00;
iconPixArray[1798] = 12'h 00;
iconPixArray[1799] = 12'h 00;
iconPixArray[1800] = 12'h 00;
iconPixArray[1801] = 12'h 00;
iconPixArray[1802] = 12'h100;
iconPixArray[1803] = 12'hE30;
iconPixArray[1804] = 12'hF30;
iconPixArray[1805] = 12'hE30;
iconPixArray[1806] = 12'hF60;
iconPixArray[1807] = 12'hE50;
iconPixArray[1808] = 12'hF60;
iconPixArray[1809] = 12'hE30;
iconPixArray[1810] = 12'hF30;
iconPixArray[1811] = 12'hB20;
iconPixArray[1812] = 12'h 00;
iconPixArray[1813] = 12'h 00;
iconPixArray[1814] = 12'h 00;
iconPixArray[1815] = 12'h 00;
iconPixArray[1816] = 12'h 00;
iconPixArray[1817] = 12'h 00;
iconPixArray[1818] = 12'h 00;
iconPixArray[1819] = 12'h 00;
iconPixArray[1820] = 12'h 00;
iconPixArray[1821] = 12'h 00;
iconPixArray[1822] = 12'h 00;
iconPixArray[1823] = 12'h 00;
iconPixArray[1824] = 12'h 00;
iconPixArray[1825] = 12'h 00;
iconPixArray[1826] = 12'h 00;
iconPixArray[1827] = 12'h 00;
iconPixArray[1828] = 12'h 00;
iconPixArray[1829] = 12'h 00;
iconPixArray[1830] = 12'h 00;
iconPixArray[1831] = 12'h 00;
iconPixArray[1832] = 12'h 00;
iconPixArray[1833] = 12'h 00;
iconPixArray[1834] = 12'h100;
iconPixArray[1835] = 12'hB20;
iconPixArray[1836] = 12'h820;
iconPixArray[1837] = 12'hF30;
iconPixArray[1838] = 12'hF30;
iconPixArray[1839] = 12'hF30;
iconPixArray[1840] = 12'hF30;
iconPixArray[1841] = 12'h820;
iconPixArray[1842] = 12'hC30;
iconPixArray[1843] = 12'hD30;
iconPixArray[1844] = 12'h 00;
iconPixArray[1845] = 12'h 00;
iconPixArray[1846] = 12'h 00;
iconPixArray[1847] = 12'h 00;
iconPixArray[1848] = 12'h 00;
iconPixArray[1849] = 12'h 00;
iconPixArray[1850] = 12'h 00;
iconPixArray[1851] = 12'h 00;
iconPixArray[1852] = 12'h 00;
iconPixArray[1853] = 12'h 00;
iconPixArray[1854] = 12'h 00;
iconPixArray[1855] = 12'h 00;
iconPixArray[1856] = 12'h 00;
iconPixArray[1857] = 12'h 00;
iconPixArray[1858] = 12'h 00;
iconPixArray[1859] = 12'h 00;
iconPixArray[1860] = 12'h 00;
iconPixArray[1861] = 12'h 00;
iconPixArray[1862] = 12'h 00;
iconPixArray[1863] = 12'h 00;
iconPixArray[1864] = 12'h 00;
iconPixArray[1865] = 12'h 00;
iconPixArray[1866] = 12'h 00;
iconPixArray[1867] = 12'h 00;
iconPixArray[1868] = 12'h410;
iconPixArray[1869] = 12'hE40;
iconPixArray[1870] = 12'hD30;
iconPixArray[1871] = 12'h920;
iconPixArray[1872] = 12'hF40;
iconPixArray[1873] = 12'h510;
iconPixArray[1874] = 12'h200;
iconPixArray[1875] = 12'h820;
iconPixArray[1876] = 12'h 00;
iconPixArray[1877] = 12'h 00;
iconPixArray[1878] = 12'h 00;
iconPixArray[1879] = 12'h 00;
iconPixArray[1880] = 12'h 00;
iconPixArray[1881] = 12'h 00;
iconPixArray[1882] = 12'h 00;
iconPixArray[1883] = 12'h 00;
iconPixArray[1884] = 12'h 00;
iconPixArray[1885] = 12'h 00;
iconPixArray[1886] = 12'h 00;
iconPixArray[1887] = 12'h 00;
iconPixArray[1888] = 12'h 00;
iconPixArray[1889] = 12'h 00;
iconPixArray[1890] = 12'h 00;
iconPixArray[1891] = 12'h 00;
iconPixArray[1892] = 12'h 00;
iconPixArray[1893] = 12'h 00;
iconPixArray[1894] = 12'h 00;
iconPixArray[1895] = 12'h 00;
iconPixArray[1896] = 12'h 00;
iconPixArray[1897] = 12'h 00;
iconPixArray[1898] = 12'h 00;
iconPixArray[1899] = 12'h 00;
iconPixArray[1900] = 12'h300;
iconPixArray[1901] = 12'hF40;
iconPixArray[1902] = 12'h920;
iconPixArray[1903] = 12'h 00;
iconPixArray[1904] = 12'hE30;
iconPixArray[1905] = 12'h610;
iconPixArray[1906] = 12'h 00;
iconPixArray[1907] = 12'h 00;
iconPixArray[1908] = 12'h 00;
iconPixArray[1909] = 12'h 00;
iconPixArray[1910] = 12'h 00;
iconPixArray[1911] = 12'h 00;
iconPixArray[1912] = 12'h 00;
iconPixArray[1913] = 12'h 00;
iconPixArray[1914] = 12'h 00;
iconPixArray[1915] = 12'h 00;
iconPixArray[1916] = 12'h 00;
iconPixArray[1917] = 12'h 00;
iconPixArray[1918] = 12'h 00;
iconPixArray[1919] = 12'h 00;
iconPixArray[1920] = 12'h 00;
iconPixArray[1921] = 12'h 00;
iconPixArray[1922] = 12'h 00;
iconPixArray[1923] = 12'h 00;
iconPixArray[1924] = 12'h 00;
iconPixArray[1925] = 12'h 00;
iconPixArray[1926] = 12'h 00;
iconPixArray[1927] = 12'h 00;
iconPixArray[1928] = 12'h 00;
iconPixArray[1929] = 12'h 00;
iconPixArray[1930] = 12'h 00;
iconPixArray[1931] = 12'h 00;
iconPixArray[1932] = 12'h100;
iconPixArray[1933] = 12'hE30;
iconPixArray[1934] = 12'h300;
iconPixArray[1935] = 12'h 00;
iconPixArray[1936] = 12'h820;
iconPixArray[1937] = 12'h510;
iconPixArray[1938] = 12'h 00;
iconPixArray[1939] = 12'h 00;
iconPixArray[1940] = 12'h 00;
iconPixArray[1941] = 12'h 00;
iconPixArray[1942] = 12'h 00;
iconPixArray[1943] = 12'h 00;
iconPixArray[1944] = 12'h 00;
iconPixArray[1945] = 12'h 00;
iconPixArray[1946] = 12'h 00;
iconPixArray[1947] = 12'h 00;
iconPixArray[1948] = 12'h 00;
iconPixArray[1949] = 12'h 00;
iconPixArray[1950] = 12'h 00;
iconPixArray[1951] = 12'h 00;
iconPixArray[1952] = 12'h 00;
iconPixArray[1953] = 12'h 00;
iconPixArray[1954] = 12'h 00;
iconPixArray[1955] = 12'h 00;
iconPixArray[1956] = 12'h 00;
iconPixArray[1957] = 12'h 00;
iconPixArray[1958] = 12'h 00;
iconPixArray[1959] = 12'h 00;
iconPixArray[1960] = 12'h 00;
iconPixArray[1961] = 12'h 00;
iconPixArray[1962] = 12'h 00;
iconPixArray[1963] = 12'h 00;
iconPixArray[1964] = 12'h 00;
iconPixArray[1965] = 12'h200;
iconPixArray[1966] = 12'h 00;
iconPixArray[1967] = 12'h 00;
iconPixArray[1968] = 12'h 00;
iconPixArray[1969] = 12'h 00;
iconPixArray[1970] = 12'h 00;
iconPixArray[1971] = 12'h 00;
iconPixArray[1972] = 12'h 00;
iconPixArray[1973] = 12'h 00;
iconPixArray[1974] = 12'h 00;
iconPixArray[1975] = 12'h 00;
iconPixArray[1976] = 12'h 00;
iconPixArray[1977] = 12'h 00;
iconPixArray[1978] = 12'h 00;
iconPixArray[1979] = 12'h 00;
iconPixArray[1980] = 12'h 00;
iconPixArray[1981] = 12'h 00;
iconPixArray[1982] = 12'h 00;
iconPixArray[1983] = 12'h 00;
iconPixArray[1984] = 12'h 00;
iconPixArray[1985] = 12'h 00;
iconPixArray[1986] = 12'h 00;
iconPixArray[1987] = 12'h 00;
iconPixArray[1988] = 12'h 00;
iconPixArray[1989] = 12'h 00;
iconPixArray[1990] = 12'h 00;
iconPixArray[1991] = 12'h 00;
iconPixArray[1992] = 12'h 00;
iconPixArray[1993] = 12'h 00;
iconPixArray[1994] = 12'h 00;
iconPixArray[1995] = 12'h 00;
iconPixArray[1996] = 12'h 00;
iconPixArray[1997] = 12'h 00;
iconPixArray[1998] = 12'h 00;
iconPixArray[1999] = 12'h 00;
iconPixArray[2000] = 12'h 00;
iconPixArray[2001] = 12'h 00;
iconPixArray[2002] = 12'h 00;
iconPixArray[2003] = 12'h 00;
iconPixArray[2004] = 12'h 00;
iconPixArray[2005] = 12'h 00;
iconPixArray[2006] = 12'h 00;
iconPixArray[2007] = 12'h 00;
iconPixArray[2008] = 12'h 00;
iconPixArray[2009] = 12'h 00;
iconPixArray[2010] = 12'h 00;
iconPixArray[2011] = 12'h 00;
iconPixArray[2012] = 12'h 00;
iconPixArray[2013] = 12'h 00;
iconPixArray[2014] = 12'h 00;
iconPixArray[2015] = 12'h 00;
iconPixArray[2016] = 12'h 00;
iconPixArray[2017] = 12'h 00;
iconPixArray[2018] = 12'h 00;
iconPixArray[2019] = 12'h 00;
iconPixArray[2020] = 12'h 00;
iconPixArray[2021] = 12'h 00;
iconPixArray[2022] = 12'h 00;
iconPixArray[2023] = 12'h 00;
iconPixArray[2024] = 12'h 00;
iconPixArray[2025] = 12'h 00;
iconPixArray[2026] = 12'h 00;
iconPixArray[2027] = 12'h 00;
iconPixArray[2028] = 12'h 00;
iconPixArray[2029] = 12'h 00;
iconPixArray[2030] = 12'h 00;
iconPixArray[2031] = 12'h 00;
iconPixArray[2032] = 12'h 00;
iconPixArray[2033] = 12'h 00;
iconPixArray[2034] = 12'h 00;
iconPixArray[2035] = 12'h 00;
iconPixArray[2036] = 12'h 00;
iconPixArray[2037] = 12'h 00;
iconPixArray[2038] = 12'h 00;
iconPixArray[2039] = 12'h 00;
iconPixArray[2040] = 12'h 00;
iconPixArray[2041] = 12'h 00;
iconPixArray[2042] = 12'h 00;
iconPixArray[2043] = 12'h 00;
iconPixArray[2044] = 12'h 00;
iconPixArray[2045] = 12'h 00;
iconPixArray[2046] = 12'h 00;
iconPixArray[2047] = 12'h 00;
*/
/**********************************************
*****  End of array template
***********************************************/



  end
endmodule 

:`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// filename:	icon.v
//
// ECE 540 Project 2: RojoBot World
//
// Jordan Fluth <jfluth@gmail.com>
// Paul Long pwl@pdx.edu
//
// 29 October 2014
//
// Description:
//
// 
//
//
//
//////////////////////////////////////////////////////////////////////////////////
module icon (
  
  ///////////////////////////////////////////////////////////////////////////
  // Port Declarations
  ///////////////////////////////////////////////////////////////////////////
  input					clk,
  input			[9:0]	pixCol,			// Current pixel getting drawn
  input			[9:0]	pixRow,
  input			[9:0]	locX,			// RoboCop's current location
  input			[9:0]	locY,			// top left corner
  input			[7:0]	botInfo,
  output	reg	[11:0]	botIcon			// 12-bit rgb color
);


  ///////////////////////////////////////////////////////////////////////////
  // Some Nice Constants
  ///////////////////////////////////////////////////////////////////////////
  localparam N  = 3'b000;				// These are the BotInfo_reg encodings
  localparam S  = 3'b100;				// for compass heading
  localparam E  = 3'b010;
  localparam W  = 3'b110;
  localparam NE = 3'b001;
  localparam SW = 3'b101;
  localparam SE = 3'b011;
  localparam NW = 3'b111;
  
  
  ///////////////////////////////////////////////////////////////////////////
  // Internal Signals
  ///////////////////////////////////////////////////////////////////////////
  reg	[3:0]	iconBitmapX, iconBitmapY;		// index into icon pixelmap ROM
  //reg	[3:0]	centeredLocX, centeredLocY;	// adjustment to center bot on line
  //wire	[3:0]	stretchLocX, stretchLocY;
  wire	[9:0]	iconLeft;			// Bounds of the icon 
  wire	[9:0]	iconRight;
  wire	[9:0]	iconTop;
  wire	[9:0]	iconBottom;
  
  wire	[11:0]	pixelColor;			// Color out from ROM
  reg	[8:0]	romAddress;		
  reg	[11:0]	iconPixArray[511:0];
 
  
  
  // These are the icon index transforms that need done in order to use
  // 2 Icons for the eight ordinal directions in which the bot can be headed
  wire	[8:0]	xformN  = {1'b0, 		iconBitmapY,		iconBitmapX }; 
  wire	[8:0]	xformS  = {1'b0, 4'd15-	iconBitmapY, 4'd15-	iconBitmapX }; 
  wire	[8:0]	xformE  = {1'b0, 4'd15-	iconBitmapX, 		iconBitmapY }; 
  wire	[8:0]	xformW  = {1'b0, 		iconBitmapX, 4'd15-	iconBitmapY }; 
  wire	[8:0]	xformNE = {1'b1, 		iconBitmapY, 		iconBitmapX };
  wire	[8:0]	xformSW = {1'b1, 4'd15-	iconBitmapY, 4'd15-	iconBitmapX };
  wire	[8:0]	xformSE = {1'b1, 4'd15-	iconBitmapX, 		iconBitmapY };
  wire	[8:0]	xformNW = {1'b1, 		iconBitmapX, 4'd15-	iconBitmapY };
  
  
  
  ///////////////////////////////////////////////////////////////////////////
  // Global Assigns
  ///////////////////////////////////////////////////////////////////////////
  // This give us an 16x16 box centered on both loc(x,y) and the line
  assign iconLeft   = locX-10'd6;
  assign iconRight  = locX+10'd9;
  assign iconTop    = locY-10'd6;
  assign iconBottom = locY+10'd9;
  
 
  ///////////////////////////////////////////////////////////////////////////
  // Instantiate the Block ROM holding Icon
  ///////////////////////////////////////////////////////////////////////////
  /*iconRom iconROM (
	.clka	(clk),
	.ena	(1'b0),				// Always enabled
	.addra	(romAddress),
	.douta	(pixelColor));*/
  
  
  // Set index into icon
  always @ (posedge clk) begin
	iconBitmapX <= pixCol[3:0] - iconLeft[3:0];
	iconBitmapY <= pixRow[3:0] -  iconTop[3:0];
  end
  
 
  // Decide when to paint the botIcon
  // If the cathode ray gun overlaps the adjusted bot location,
  // paint the icon, otherwise paint "00" (transparency)

  always @ (posedge clk) begin
	if (pixCol >= iconLeft && pixCol <= iconRight &&
		pixRow >= iconTop  && pixRow <= iconBottom) begin
		
		case (botInfo[2:0])
			N :	botIcon <= iconPixArray[xformN];
			S :	botIcon <= iconPixArray[xformS];
			E :	botIcon <= iconPixArray[xformE];
			W :	botIcon <= iconPixArray[xformW];
			NE:	botIcon <= iconPixArray[xformNE];
			NW:	botIcon <= iconPixArray[xformNW];
			SE:	botIcon <= iconPixArray[xformSE];
			SW:	botIcon <= iconPixArray[xformSW];
			// We should never get here
			default: botIcon <= 12'b0;
		endcase	
	end
	else begin
		botIcon    <= 12'b0;				// transparent 
	end
  end
	  
  initial begin
                          

	/*
	// Block Arrow
	iconPixArray[0]   = 12'hf00;
	iconPixArray[1]   = 12'hf00;
	iconPixArray[2]   = 12'hf00;
	iconPixArray[3]   = 12'hf00;
	iconPixArray[4]   = 12'hf00;
	iconPixArray[5]   = 12'hf00;
	iconPixArray[6]   = 12'hf00;
	iconPixArray[7]   = 12'hf00;
	iconPixArray[8]   = 12'hf00;
	iconPixArray[9]   = 12'hf00;
	iconPixArray[10]  = 12'hf00;
	iconPixArray[11]  = 12'hf00;
	iconPixArray[12]  = 12'hf00;
	iconPixArray[13]  = 12'hf00;
	iconPixArray[14]  = 12'hf00;
	iconPixArray[15]  = 12'hf00;
	iconPixArray[16]  = 12'hf00;
	iconPixArray[17]  = 12'hf00;
	iconPixArray[18]  = 12'hf00;
	iconPixArray[19]  = 12'hf00;
	iconPixArray[20]  = 12'hf00;
	iconPixArray[21]  = 12'hf00;
	iconPixArray[22]  = 12'hf00;
	iconPixArray[23]  = 12'hf0f;
	iconPixArray[24]  = 12'hf0f;
	iconPixArray[25]  = 12'hf00;
	iconPixArray[26]  = 12'hf00;
	iconPixArray[27]  = 12'hf00;
	iconPixArray[28]  = 12'hf00;
	iconPixArray[29]  = 12'hf00;
	iconPixArray[30]  = 12'hf00;
	iconPixArray[31]  = 12'hf00;
	iconPixArray[32]  = 12'hf00;
	iconPixArray[33]  = 12'hf00;
	iconPixArray[34]  = 12'hf00;
	iconPixArray[35]  = 12'hf00;
	iconPixArray[36]  = 12'hf00;
	iconPixArray[37]  = 12'hf00;
	iconPixArray[38]  = 12'hf0f;
	iconPixArray[39]  = 12'hf0f;
	iconPixArray[40]  = 12'hf0f;
	iconPixArray[41]  = 12'hf0f;
	iconPixArray[42]  = 12'hf00;
	iconPixArray[43]  = 12'hf00;
	iconPixArray[44]  = 12'hf00;
	iconPixArray[45]  = 12'hf00;
	iconPixArray[46]  = 12'hf00;
	iconPixArray[47]  = 12'hf00;
	iconPixArray[48]  = 12'hf00;
	iconPixArray[49]  = 12'hf00;
	iconPixArray[50]  = 12'hf00;
	iconPixArray[51]  = 12'hf00;
	iconPixArray[52]  = 12'hf00;
	iconPixArray[53]  = 12'hf0f;
	iconPixArray[54]  = 12'hf0f;
	iconPixArray[55]  = 12'hf0f;
	iconPixArray[56]  = 12'hf0f;
	iconPixArray[57]  = 12'hf0f;
	iconPixArray[58]  = 12'hf0f;
	iconPixArray[59]  = 12'hf00;
	iconPixArray[60]  = 12'hf00;
	iconPixArray[61]  = 12'hf00;
	iconPixArray[62]  = 12'hf00;
	iconPixArray[63]  = 12'hf00;
	iconPixArray[64]  = 12'hf00;
	iconPixArray[65]  = 12'hf00;
	iconPixArray[66]  = 12'hf00;
	iconPixArray[67]  = 12'hf00;
	iconPixArray[68]  = 12'hf0f;
	iconPixArray[69]  = 12'hf0f;
	iconPixArray[70]  = 12'hf0f;
	iconPixArray[71]  = 12'hf0f;
	iconPixArray[72]  = 12'hf0f;
	iconPixArray[73]  = 12'hf0f;
	iconPixArray[74]  = 12'hf0f;
	iconPixArray[75]  = 12'hf0f;
	iconPixArray[76]  = 12'hf00;
	iconPixArray[77]  = 12'hf00;
	iconPixArray[78]  = 12'hf00;
	iconPixArray[79]  = 12'hf00;
	iconPixArray[80]  = 12'hf00;
	iconPixArray[81]  = 12'hf00;
	iconPixArray[82]  = 12'hf00;
	iconPixArray[83]  = 12'hf0f;
	iconPixArray[84]  = 12'hf0f;
	iconPixArray[85]  = 12'hf0f;
	iconPixArray[86]  = 12'hf0f;
	iconPixArray[87]  = 12'hf0f;
	iconPixArray[88]  = 12'hf0f;
	iconPixArray[89]  = 12'hf0f;
	iconPixArray[90]  = 12'hf0f;
	iconPixArray[91]  = 12'hf0f;
	iconPixArray[92]  = 12'hf0f;
	iconPixArray[93]  = 12'hf00;
	iconPixArray[94]  = 12'hf00;
	iconPixArray[95]  = 12'hf00;
	iconPixArray[96]  = 12'hf00;
	iconPixArray[97]  = 12'hf00;
	iconPixArray[98]  = 12'hf0f;
	iconPixArray[99]  = 12'hf0f;
	iconPixArray[100] = 12'hf0f;
	iconPixArray[101] = 12'hf0f;
	iconPixArray[102] = 12'hf0f;
	iconPixArray[103] = 12'hf0f;
	iconPixArray[104] = 12'hf0f;
	iconPixArray[105] = 12'hf0f;
	iconPixArray[106] = 12'hf0f;
	iconPixArray[107] = 12'hf0f;
	iconPixArray[108] = 12'hf0f;
	iconPixArray[109] = 12'hf0f;
	iconPixArray[110] = 12'hf00;
	iconPixArray[111] = 12'hf00;
	iconPixArray[112] = 12'hf00;
	iconPixArray[113] = 12'hf0f;
	iconPixArray[114] = 12'hf0f;
	iconPixArray[115] = 12'hf0f;
	iconPixArray[116] = 12'hf0f;
	iconPixArray[117] = 12'hf0f;
	iconPixArray[118] = 12'hf0f;
	iconPixArray[119] = 12'hf0f;
	iconPixArray[120] = 12'hf0f;
	iconPixArray[121] = 12'hf0f;
	iconPixArray[122] = 12'hf0f;
	iconPixArray[123] = 12'hf0f;
	iconPixArray[124] = 12'hf0f;
	iconPixArray[125] = 12'hf0f;
	iconPixArray[126] = 12'hf0f;
	iconPixArray[127] = 12'hf00;
	iconPixArray[128] = 12'hf00;
	iconPixArray[129] = 12'hf00;
	iconPixArray[130] = 12'hf00;
	iconPixArray[131] = 12'hf00;
	iconPixArray[132] = 12'hf00;
	iconPixArray[133] = 12'hf0f;
	iconPixArray[134] = 12'hf0f;
	iconPixArray[135] = 12'hf0f;
	iconPixArray[136] = 12'hf0f;
	iconPixArray[137] = 12'hf0f;
	iconPixArray[138] = 12'hf0f;
	iconPixArray[139] = 12'hf00;
	iconPixArray[140] = 12'hf00;
	iconPixArray[141] = 12'hf00;
	iconPixArray[142] = 12'hf00;
	iconPixArray[143] = 12'hf00;
	iconPixArray[144] = 12'hf00;
	iconPixArray[145] = 12'hf00;
	iconPixArray[146] = 12'hf00;
	iconPixArray[147] = 12'hf00;
	iconPixArray[148] = 12'hf00;
	iconPixArray[149] = 12'hf0f;
	iconPixArray[150] = 12'hf0f;
	iconPixArray[151] = 12'hf0f;
	iconPixArray[152] = 12'hf0f;
	iconPixArray[153] = 12'hf0f;
	iconPixArray[154] = 12'hf0f;
	iconPixArray[155] = 12'hf00;
	iconPixArray[156] = 12'hf00;
	iconPixArray[157] = 12'hf00;
	iconPixArray[158] = 12'hf00;
	iconPixArray[159] = 12'hf00;
	iconPixArray[160] = 12'hf00;
	iconPixArray[161] = 12'hf00;
	iconPixArray[162] = 12'hf00;
	iconPixArray[163] = 12'hf00;
	iconPixArray[164] = 12'hf00;
	iconPixArray[165] = 12'hf0f;
	iconPixArray[166] = 12'hf0f;
	iconPixArray[167] = 12'hf0f;
	iconPixArray[168] = 12'hf0f;
	iconPixArray[169] = 12'hf0f;
	iconPixArray[170] = 12'hf0f;
	iconPixArray[171] = 12'hf00;
	iconPixArray[172] = 12'hf00;
	iconPixArray[173] = 12'hf00;
	iconPixArray[174] = 12'hf00;
	iconPixArray[175] = 12'hf00;
	iconPixArray[176] = 12'hf00;
	iconPixArray[177] = 12'hf00;
	iconPixArray[178] = 12'hf00;
	iconPixArray[179] = 12'hf00;
	iconPixArray[180] = 12'hf00;
	iconPixArray[181] = 12'hf0f;
	iconPixArray[182] = 12'hf0f;
	iconPixArray[183] = 12'hf0f;
	iconPixArray[184] = 12'hf0f;
	iconPixArray[185] = 12'hf0f;
	iconPixArray[186] = 12'hf0f;
	iconPixArray[187] = 12'hf00;
	iconPixArray[188] = 12'hf00;
	iconPixArray[189] = 12'hf00;
	iconPixArray[190] = 12'hf00;
	iconPixArray[191] = 12'hf00;
	iconPixArray[192] = 12'hf00;
	iconPixArray[193] = 12'hf00;
	iconPixArray[194] = 12'hf00;
	iconPixArray[195] = 12'hf00;
	iconPixArray[196] = 12'hf00;
	iconPixArray[197] = 12'hf0f;
	iconPixArray[198] = 12'hf0f;
	iconPixArray[199] = 12'hf0f;
	iconPixArray[200] = 12'hf0f;
	iconPixArray[201] = 12'hf0f;
	iconPixArray[202] = 12'hf0f;
	iconPixArray[203] = 12'hf00;
	iconPixArray[204] = 12'hf00;
	iconPixArray[205] = 12'hf00;
	iconPixArray[206] = 12'hf00;
	iconPixArray[207] = 12'hf00;
	iconPixArray[208] = 12'hf00;
	iconPixArray[209] = 12'hf00;
	iconPixArray[210] = 12'hf00;
	iconPixArray[211] = 12'hf00;
	iconPixArray[212] = 12'hf00;
	iconPixArray[213] = 12'hf0f;
	iconPixArray[214] = 12'hf0f;
	iconPixArray[215] = 12'hf0f;
	iconPixArray[216] = 12'hf0f;
	iconPixArray[217] = 12'hf0f;
	iconPixArray[218] = 12'hf0f;
	iconPixArray[219] = 12'hf00;
	iconPixArray[220] = 12'hf00;
	iconPixArray[221] = 12'hf00;
	iconPixArray[222] = 12'hf00;
	iconPixArray[223] = 12'hf00;
	iconPixArray[224] = 12'hf00;
	iconPixArray[225] = 12'hf00;
	iconPixArray[226] = 12'hf00;
	iconPixArray[227] = 12'hf00;
	iconPixArray[228] = 12'hf00;
	iconPixArray[229] = 12'hf0f;
	iconPixArray[230] = 12'hf0f;
	iconPixArray[231] = 12'hf0f;
	iconPixArray[232] = 12'hf0f;
	iconPixArray[233] = 12'hf0f;
	iconPixArray[234] = 12'hf0f;
	iconPixArray[235] = 12'hf00;
	iconPixArray[236] = 12'hf00;
	iconPixArray[237] = 12'hf00;
	iconPixArray[238] = 12'hf00;
	iconPixArray[239] = 12'hf00;
	iconPixArray[240] = 12'hf00;
	iconPixArray[241] = 12'hf00;
	iconPixArray[242] = 12'hf00;
	iconPixArray[243] = 12'hf00;
	iconPixArray[244] = 12'hf00;
	iconPixArray[245] = 12'hf00;
	iconPixArray[246] = 12'hf00;
	iconPixArray[247] = 12'hf00;
	iconPixArray[248] = 12'hf00;
	iconPixArray[249] = 12'hf00;
	iconPixArray[250] = 12'hf00;
	iconPixArray[251] = 12'hf00;
	iconPixArray[252] = 12'hf00;
	iconPixArray[253] = 12'hf00;
	iconPixArray[254] = 12'hf00;
	iconPixArray[255] = 12'hf00;	

	iconPixArray[256] = 12'hf00;
	iconPixArray[257] = 12'hf00;
	iconPixArray[258] = 12'hf00;
	iconPixArray[259] = 12'hf00;
	iconPixArray[260] = 12'hf00;
	iconPixArray[261] = 12'hf00;
	iconPixArray[262] = 12'hf00;
	iconPixArray[263] = 12'hf00;
	iconPixArray[264] = 12'hf00;
	iconPixArray[265] = 12'hf00;
	iconPixArray[266] = 12'hf00;
	iconPixArray[267] = 12'hf00;
	iconPixArray[268] = 12'hf00;
	iconPixArray[269] = 12'hf00;
	iconPixArray[270] = 12'hf00;
	iconPixArray[271] = 12'hf00;
	iconPixArray[272] = 12'hf00;
	iconPixArray[273] = 12'hf00;
	iconPixArray[274] = 12'hf00;
	iconPixArray[275] = 12'hf0f;
	iconPixArray[276] = 12'hf0f;
	iconPixArray[277] = 12'hf0f;
	iconPixArray[278] = 12'hf0f;
	iconPixArray[279] = 12'hf0f;
	iconPixArray[280] = 12'hf0f;
	iconPixArray[281] = 12'hf0f;
	iconPixArray[282] = 12'hf0f;
	iconPixArray[283] = 12'hf0f;
	iconPixArray[284] = 12'hf0f;
	iconPixArray[285] = 12'hf0f;
	iconPixArray[286] = 12'hf0f;
	iconPixArray[287] = 12'hf00;
	iconPixArray[288] = 12'hf00;
	iconPixArray[289] = 12'hf00;
	iconPixArray[290] = 12'hf00;
	iconPixArray[291] = 12'hf00;
	iconPixArray[292] = 12'hf00;
	iconPixArray[293] = 12'hf0f;
	iconPixArray[294] = 12'hf0f;
	iconPixArray[295] = 12'hf0f;
	iconPixArray[296] = 12'hf0f;
	iconPixArray[297] = 12'hf0f;
	iconPixArray[298] = 12'hf0f;
	iconPixArray[299] = 12'hf0f;
	iconPixArray[300] = 12'hf0f;
	iconPixArray[301] = 12'hf0f;
	iconPixArray[302] = 12'hf0f;
	iconPixArray[303] = 12'hf00;
	iconPixArray[304] = 12'hf00;
	iconPixArray[305] = 12'hf00;
	iconPixArray[306] = 12'hf00;
	iconPixArray[307] = 12'hf00;
	iconPixArray[308] = 12'hf00;
	iconPixArray[309] = 12'hf00;
	iconPixArray[310] = 12'hf00;
	iconPixArray[311] = 12'hf0f;
	iconPixArray[312] = 12'hf0f;
	iconPixArray[313] = 12'hf0f;
	iconPixArray[314] = 12'hf0f;
	iconPixArray[315] = 12'hf0f;
	iconPixArray[316] = 12'hf0f;
	iconPixArray[317] = 12'hf0f;
	iconPixArray[318] = 12'hf0f;
	iconPixArray[319] = 12'hf00;
	iconPixArray[320] = 12'hf00;
	iconPixArray[321] = 12'hf00;
	iconPixArray[322] = 12'hf00;
	iconPixArray[323] = 12'hf00;
	iconPixArray[324] = 12'hf00;
	iconPixArray[325] = 12'hf00;
	iconPixArray[326] = 12'hf00;
	iconPixArray[327] = 12'hf00;
	iconPixArray[328] = 12'hf00;
	iconPixArray[329] = 12'hf0f;
	iconPixArray[330] = 12'hf0f;
	iconPixArray[331] = 12'hf0f;
	iconPixArray[332] = 12'hf0f;
	iconPixArray[333] = 12'hf0f;
	iconPixArray[334] = 12'hf0f;
	iconPixArray[335] = 12'hf00;
	iconPixArray[336] = 12'hf00;
	iconPixArray[337] = 12'hf00;
	iconPixArray[338] = 12'hf00;
	iconPixArray[339] = 12'hf00;
	iconPixArray[340] = 12'hf00;
	iconPixArray[341] = 12'hf00;
	iconPixArray[342] = 12'hf00;
	iconPixArray[343] = 12'hf00;
	iconPixArray[344] = 12'hf00;
	iconPixArray[345] = 12'hf0f;
	iconPixArray[346] = 12'hf0f;
	iconPixArray[347] = 12'hf0f;
	iconPixArray[348] = 12'hf0f;
	iconPixArray[349] = 12'hf0f;
	iconPixArray[350] = 12'hf0f;
	iconPixArray[351] = 12'hf00;
	iconPixArray[352] = 12'hf00;
	iconPixArray[353] = 12'hf00;
	iconPixArray[354] = 12'hf00;
	iconPixArray[355] = 12'hf00;
	iconPixArray[356] = 12'hf00;
	iconPixArray[357] = 12'hf00;
	iconPixArray[358] = 12'hf00;
	iconPixArray[359] = 12'hf00;
	iconPixArray[360] = 12'hf0f;
	iconPixArray[361] = 12'hf0f;
	iconPixArray[362] = 12'hf0f;
	iconPixArray[363] = 12'hf0f;
	iconPixArray[364] = 12'hf0f;
	iconPixArray[365] = 12'hf0f;
	iconPixArray[366] = 12'hf0f;
	iconPixArray[367] = 12'hf00;
	iconPixArray[368] = 12'hf00;
	iconPixArray[369] = 12'hf00;
	iconPixArray[370] = 12'hf00;
	iconPixArray[371] = 12'hf00;
	iconPixArray[372] = 12'hf00;
	iconPixArray[373] = 12'hf00;
	iconPixArray[374] = 12'hf00;
	iconPixArray[375] = 12'hf0f;
	iconPixArray[376] = 12'hf0f;
	iconPixArray[377] = 12'hf0f;
	iconPixArray[378] = 12'hf00;
	iconPixArray[379] = 12'hf00;
	iconPixArray[380] = 12'hf0f;
	iconPixArray[381] = 12'hf0f;
	iconPixArray[382] = 12'hf0f;
	iconPixArray[383] = 12'hf00;
	iconPixArray[384] = 12'hf00;
	iconPixArray[385] = 12'hf00;
	iconPixArray[386] = 12'hf00;
	iconPixArray[387] = 12'hf00;
	iconPixArray[388] = 12'hf00;
	iconPixArray[389] = 12'hf00;
	iconPixArray[390] = 12'hf0f;
	iconPixArray[391] = 12'hf0f;
	iconPixArray[392] = 12'hf0f;
	iconPixArray[393] = 12'hf00;
	iconPixArray[394] = 12'hf00;
	iconPixArray[395] = 12'hf00;
	iconPixArray[396] = 12'hf0f;
	iconPixArray[397] = 12'hf0f;
	iconPixArray[398] = 12'hf0f;
	iconPixArray[399] = 12'hf00;
	iconPixArray[400] = 12'hf00;
	iconPixArray[401] = 12'hf00;
	iconPixArray[402] = 12'hf00;
	iconPixArray[403] = 12'hf00;
	iconPixArray[404] = 12'hf00;
	iconPixArray[405] = 12'hf0f;
	iconPixArray[406] = 12'hf0f;
	iconPixArray[407] = 12'hf0f;
	iconPixArray[408] = 12'hf00;
	iconPixArray[409] = 12'hf00;
	iconPixArray[410] = 12'hf00;
	iconPixArray[411] = 12'hf00;
	iconPixArray[412] = 12'hf0f;
	iconPixArray[413] = 12'hf0f;
	iconPixArray[414] = 12'hf0f;
	iconPixArray[415] = 12'hf00;
	iconPixArray[416] = 12'hf00;
	iconPixArray[417] = 12'hf00;
	iconPixArray[418] = 12'hf00;
	iconPixArray[419] = 12'hf00;
	iconPixArray[420] = 12'hf0f;
	iconPixArray[421] = 12'hf0f;
	iconPixArray[422] = 12'hf0f;
	iconPixArray[423] = 12'hf00;
	iconPixArray[424] = 12'hf00;
	iconPixArray[425] = 12'hf00;
	iconPixArray[426] = 12'hf00;
	iconPixArray[427] = 12'hf00;
	iconPixArray[428] = 12'hf00;
	iconPixArray[429] = 12'hf0f;
	iconPixArray[430] = 12'hf0f;
	iconPixArray[431] = 12'hf00;
	iconPixArray[432] = 12'hf00;
	iconPixArray[433] = 12'hf00;
	iconPixArray[434] = 12'hf00;
	iconPixArray[435] = 12'hf0f;
	iconPixArray[436] = 12'hf0f;
	iconPixArray[437] = 12'hf00;
	iconPixArray[438] = 12'hf00;
	iconPixArray[439] = 12'hf00;
	iconPixArray[440] = 12'hf00;
	iconPixArray[441] = 12'hf00;
	iconPixArray[442] = 12'hf00;
	iconPixArray[443] = 12'hf00;
	iconPixArray[444] = 12'hf00;
	iconPixArray[445] = 12'hf00;
	iconPixArray[446] = 12'hf0f;
	iconPixArray[447] = 12'hf00;
	iconPixArray[448] = 12'hf00;
	iconPixArray[449] = 12'hf00;
	iconPixArray[450] = 12'hf0f;
	iconPixArray[451] = 12'hf0f;
	iconPixArray[452] = 12'hf0f;
	iconPixArray[453] = 12'hf00;
	iconPixArray[454] = 12'hf00;
	iconPixArray[455] = 12'hf00;
	iconPixArray[456] = 12'hf00;
	iconPixArray[457] = 12'hf00;
	iconPixArray[458] = 12'hf00;
	iconPixArray[459] = 12'hf00;
	iconPixArray[460] = 12'hf00;
	iconPixArray[461] = 12'hf00;
	iconPixArray[462] = 12'hf0f;
	iconPixArray[463] = 12'hf00;
	iconPixArray[464] = 12'hf00;
	iconPixArray[465] = 12'hf0f;
	iconPixArray[466] = 12'hf0f;
	iconPixArray[467] = 12'hf0f;
	iconPixArray[468] = 12'hf00;
	iconPixArray[469] = 12'hf00;
	iconPixArray[470] = 12'hf00;
	iconPixArray[471] = 12'hf00;
	iconPixArray[472] = 12'hf00;
	iconPixArray[473] = 12'hf00;
	iconPixArray[474] = 12'hf00;
	iconPixArray[475] = 12'hf00;
	iconPixArray[476] = 12'hf00;
	iconPixArray[477] = 12'hf00;
	iconPixArray[478] = 12'hf00;
	iconPixArray[479] = 12'hf00;
	iconPixArray[480] = 12'hf00;
	iconPixArray[481] = 12'hf0f;
	iconPixArray[482] = 12'hf0f;
	iconPixArray[483] = 12'hf00;
	iconPixArray[484] = 12'hf00;
	iconPixArray[485] = 12'hf00;
	iconPixArray[486] = 12'hf00;
	iconPixArray[487] = 12'hf00;
	iconPixArray[488] = 12'hf00;
	iconPixArray[489] = 12'hf00;
	iconPixArray[490] = 12'hf00;
	iconPixArray[491] = 12'hf00;
	iconPixArray[492] = 12'hf00;
	iconPixArray[493] = 12'hf00;
	iconPixArray[494] = 12'hf00;
	iconPixArray[495] = 12'hf00;
	iconPixArray[496] = 12'hf00;
	iconPixArray[497] = 12'hf00;
	iconPixArray[498] = 12'hf00;
	iconPixArray[499] = 12'hf00;
	iconPixArray[500] = 12'hf00;
	iconPixArray[501] = 12'hf00;
	iconPixArray[502] = 12'hf00;
	iconPixArray[503] = 12'hf00;
	iconPixArray[504] = 12'hf00;
	iconPixArray[505] = 12'hf00;
	iconPixArray[506] = 12'hf00;
	iconPixArray[507] = 12'hf00;
	iconPixArray[508] = 12'hf00;
	iconPixArray[509] = 12'hf00;
	iconPixArray[510] = 12'hf00;
	iconPixArray[511] = 12'hf00;
<<<<<<< HEAD
 */                 
                 


/*
//skull
iconPixArray[0] = 12'h000;
iconPixArray[1] = 12'h000;
iconPixArray[2] = 12'h000;
iconPixArray[3] = 12'h000;
iconPixArray[4] = 12'h000;
iconPixArray[5] = 12'h5BB;
iconPixArray[6] = 12'h5BB;
iconPixArray[7] = 12'h5BB;
iconPixArray[8] = 12'h5BB;
iconPixArray[9] = 12'h5BB;
iconPixArray[10] = 12'h5BB;
iconPixArray[11] = 12'h000;
iconPixArray[12] = 12'h000;
iconPixArray[13] = 12'h000;
iconPixArray[14] = 12'h000;
iconPixArray[15] = 12'h000;
iconPixArray[16] = 12'h000;
iconPixArray[17] = 12'h000;
iconPixArray[18] = 12'h000;
iconPixArray[19] = 12'h5BB;
iconPixArray[20] = 12'h5BB;
iconPixArray[21] = 12'h6AA;
iconPixArray[22] = 12'hE22;
iconPixArray[23] = 12'hECC;
iconPixArray[24] = 12'hECC;
iconPixArray[25] = 12'hE22;
iconPixArray[26] = 12'h6AA;
iconPixArray[27] = 12'h5BB;
iconPixArray[28] = 12'h5BB;
iconPixArray[29] = 12'h000;
iconPixArray[30] = 12'h000;
iconPixArray[31] = 12'h000;
iconPixArray[32] = 12'h000;
iconPixArray[33] = 12'h000;
iconPixArray[34] = 12'h5BB;
iconPixArray[35] = 12'h5AA;
iconPixArray[36] = 12'hD44;
iconPixArray[37] = 12'hC00;
iconPixArray[38] = 12'hC77;
iconPixArray[39] = 12'hC33;
iconPixArray[40] = 12'hC33;
iconPixArray[41] = 12'hC77;
iconPixArray[42] = 12'hC00;
iconPixArray[43] = 12'hD44;
iconPixArray[44] = 12'h5AA;
iconPixArray[45] = 12'h5BB;
iconPixArray[46] = 12'h000;
iconPixArray[47] = 12'h000;
iconPixArray[48] = 12'h000;
iconPixArray[49] = 12'h5BB;
iconPixArray[50] = 12'h588;
iconPixArray[51] = 12'hB44;
iconPixArray[52] = 12'hAFF;
iconPixArray[53] = 12'h933;
iconPixArray[54] = 12'h9FF;
iconPixArray[55] = 12'h9FF;
iconPixArray[56] = 12'h9FF;
iconPixArray[57] = 12'h9FF;
iconPixArray[58] = 12'h9FF;
iconPixArray[59] = 12'h988;
iconPixArray[60] = 12'hB00;
iconPixArray[61] = 12'h588;
iconPixArray[62] = 12'h5BB;
iconPixArray[63] = 12'h000;
iconPixArray[64] = 12'h000;
iconPixArray[65] = 12'h5BB;
iconPixArray[66] = 12'h9BB;
iconPixArray[67] = 12'h6AA;
iconPixArray[68] = 12'h477;
iconPixArray[69] = 12'hFFF;
iconPixArray[70] = 12'hFFF;
iconPixArray[71] = 12'hFFF;
iconPixArray[72] = 12'hFFF;
iconPixArray[73] = 12'hFFF;
iconPixArray[74] = 12'hFFF;
iconPixArray[75] = 12'hFFF;
iconPixArray[76] = 12'h4BB;
iconPixArray[77] = 12'h977;
iconPixArray[78] = 12'h5BB;
iconPixArray[79] = 12'h000;
iconPixArray[80] = 12'h5BB;
iconPixArray[81] = 12'h433;
iconPixArray[82] = 12'h511;
iconPixArray[83] = 12'h288;
iconPixArray[84] = 12'hFFF;
iconPixArray[85] = 12'hFFF;
iconPixArray[86] = 12'hFFF;
iconPixArray[87] = 12'hFFF;
iconPixArray[88] = 12'hFFF;
iconPixArray[89] = 12'hFFF;
iconPixArray[90] = 12'hFFF;
iconPixArray[91] = 12'hFFF;
iconPixArray[92] = 12'hFFF;
iconPixArray[93] = 12'h366;
iconPixArray[94] = 12'h433;
iconPixArray[95] = 12'h5BB;
iconPixArray[96] = 12'h5BB;
iconPixArray[97] = 12'h6BB;
iconPixArray[98] = 12'h222;
iconPixArray[99] = 12'hFFF;
iconPixArray[100] = 12'hFFF;
iconPixArray[101] = 12'hD55;
iconPixArray[102] = 12'hD55;
iconPixArray[103] = 12'hFFF;
iconPixArray[104] = 12'hFFF;
iconPixArray[105] = 12'hFFF;
iconPixArray[106] = 12'hD55;
iconPixArray[107] = 12'hD55;
iconPixArray[108] = 12'hFFF;
iconPixArray[109] = 12'hF44;
iconPixArray[110] = 12'h6BB;
iconPixArray[111] = 12'h5BB;
iconPixArray[112] = 12'h5BB;
iconPixArray[113] = 12'h4EE;
iconPixArray[114] = 12'hF66;
iconPixArray[115] = 12'hB99;
iconPixArray[116] = 12'hFFF;
iconPixArray[117] = 12'h800;
iconPixArray[118] = 12'h800;
iconPixArray[119] = 12'hFFF;
iconPixArray[120] = 12'hFFF;
iconPixArray[121] = 12'hFFF;
iconPixArray[122] = 12'h800;
iconPixArray[123] = 12'h800;
iconPixArray[124] = 12'hFFF;
iconPixArray[125] = 12'hB99;
iconPixArray[126] = 12'h4EE;
iconPixArray[127] = 12'h5BB;
iconPixArray[128] = 12'h5BB;
iconPixArray[129] = 12'h188;
iconPixArray[130] = 12'hB00;
iconPixArray[131] = 12'h644;
iconPixArray[132] = 12'hFFF;
iconPixArray[133] = 12'hFFF;
iconPixArray[134] = 12'hFFF;
iconPixArray[135] = 12'hFFF;
iconPixArray[136] = 12'hFFF;
iconPixArray[137] = 12'hFFF;
iconPixArray[138] = 12'hFFF;
iconPixArray[139] = 12'hFFF;
iconPixArray[140] = 12'hFFF;
iconPixArray[141] = 12'h644;
iconPixArray[142] = 12'h188;
iconPixArray[143] = 12'h5BB;
iconPixArray[144] = 12'h5BB;
iconPixArray[145] = 12'h088;
iconPixArray[146] = 12'h9EE;
iconPixArray[147] = 12'h411;
iconPixArray[148] = 12'hFFF;
iconPixArray[149] = 12'hFFF;
iconPixArray[150] = 12'hFFF;
iconPixArray[151] = 12'hFFF;
iconPixArray[152] = 12'hD22;
iconPixArray[153] = 12'hFFF;
iconPixArray[154] = 12'hFFF;
iconPixArray[155] = 12'hFFF;
iconPixArray[156] = 12'hFFF;
iconPixArray[157] = 12'h555;
iconPixArray[158] = 12'h088;
iconPixArray[159] = 12'h5BB;
iconPixArray[160] = 12'h5BB;
iconPixArray[161] = 12'h166;
iconPixArray[162] = 12'h811;
iconPixArray[163] = 12'h400;
iconPixArray[164] = 12'hE66;
iconPixArray[165] = 12'hFFF;
iconPixArray[166] = 12'hFFF;
iconPixArray[167] = 12'hFFF;
iconPixArray[168] = 12'hFFF;
iconPixArray[169] = 12'hFFF;
iconPixArray[170] = 12'hFFF;
iconPixArray[171] = 12'hFFF;
iconPixArray[172] = 12'hE66;
iconPixArray[173] = 12'h7EE;
iconPixArray[174] = 12'h166;
iconPixArray[175] = 12'h5BB;
iconPixArray[176] = 12'h000;
iconPixArray[177] = 12'h5BB;
iconPixArray[178] = 12'hB00;
iconPixArray[179] = 12'h422;
iconPixArray[180] = 12'h1BB;
iconPixArray[181] = 12'hAFF;
iconPixArray[182] = 12'hFFF;
iconPixArray[183] = 12'h6AA;
iconPixArray[184] = 12'hFFF;
iconPixArray[185] = 12'h6AA;
iconPixArray[186] = 12'hFFF;
iconPixArray[187] = 12'hAFF;
iconPixArray[188] = 12'h2FF;
iconPixArray[189] = 12'hB00;
iconPixArray[190] = 12'h5BB;
iconPixArray[191] = 12'h000;
iconPixArray[192] = 12'h000;
iconPixArray[193] = 12'h5BB;
iconPixArray[194] = 12'hF11;
iconPixArray[195] = 12'h5DD;
iconPixArray[196] = 12'h1BB;
iconPixArray[197] = 12'hB11;
iconPixArray[198] = 12'hFFF;
iconPixArray[199] = 12'h6AA;
iconPixArray[200] = 12'hFFF;
iconPixArray[201] = 12'h6AA;
iconPixArray[202] = 12'hFFF;
iconPixArray[203] = 12'hC44;
iconPixArray[204] = 12'h5DD;
iconPixArray[205] = 12'hF11;
iconPixArray[206] = 12'h5BB;
iconPixArray[207] = 12'h000;
iconPixArray[208] = 12'h000;
iconPixArray[209] = 12'h000;
iconPixArray[210] = 12'h5BB;
iconPixArray[211] = 12'hEEE;
iconPixArray[212] = 12'h622;
iconPixArray[213] = 12'hFDD;
iconPixArray[214] = 12'hA22;
iconPixArray[215] = 12'h9EE;
iconPixArray[216] = 12'h9EE;
iconPixArray[217] = 12'hA22;
iconPixArray[218] = 12'hEAA;
iconPixArray[219] = 12'h5FF;
iconPixArray[220] = 12'hEEE;
iconPixArray[221] = 12'h5BB;
iconPixArray[222] = 12'h000;
iconPixArray[223] = 12'h000;
iconPixArray[224] = 12'h000;
iconPixArray[225] = 12'h000;
iconPixArray[226] = 12'h000;
iconPixArray[227] = 12'h5BB;
iconPixArray[228] = 12'h5BB;
iconPixArray[229] = 12'hE99;
iconPixArray[230] = 12'h744;
iconPixArray[231] = 12'h6EE;
iconPixArray[232] = 12'h6EE;
iconPixArray[233] = 12'h744;
iconPixArray[234] = 12'hE99;
iconPixArray[235] = 12'h5BB;
iconPixArray[236] = 12'h5BB;
iconPixArray[237] = 12'h000;
iconPixArray[238] = 12'h000;
iconPixArray[239] = 12'h000;
iconPixArray[240] = 12'h000;
iconPixArray[241] = 12'h000;
iconPixArray[242] = 12'h000;
iconPixArray[243] = 12'h000;
iconPixArray[244] = 12'h000;
iconPixArray[245] = 12'h5BB;
iconPixArray[246] = 12'h5BB;
iconPixArray[247] = 12'h5BB;
iconPixArray[248] = 12'h5BB;
iconPixArray[249] = 12'h5BB;
iconPixArray[250] = 12'h5BB;
iconPixArray[251] = 12'h000;
iconPixArray[252] = 12'h000;
iconPixArray[253] = 12'h000;
iconPixArray[254] = 12'h000;
iconPixArray[255] = 12'h000;
*/

/**********************************************
*****  Template file for the image array
*****  Produced from rocket.png
***********************************************/
/*
iconPixArray[0] = 12'h000;
iconPixArray[1] = 12'h000;
iconPixArray[2] = 12'h000;
iconPixArray[3] = 12'h000;
iconPixArray[4] = 12'h000;
iconPixArray[5] = 12'h000;
iconPixArray[6] = 12'h000;
iconPixArray[7] = 12'h000;
iconPixArray[8] = 12'h000;
iconPixArray[9] = 12'h000;
iconPixArray[10] = 12'h000;
iconPixArray[11] = 12'h000;
iconPixArray[12] = 12'h000;
iconPixArray[13] = 12'h000;
iconPixArray[14] = 12'h000;
iconPixArray[15] = 12'h000;
iconPixArray[16] = 12'h000;
iconPixArray[17] = 12'h000;
iconPixArray[18] = 12'h000;
iconPixArray[19] = 12'h000;
iconPixArray[20] = 12'h000;
iconPixArray[21] = 12'h000;
iconPixArray[22] = 12'h000;
iconPixArray[23] = 12'h000;
iconPixArray[24] = 12'h000;
iconPixArray[25] = 12'h000;
iconPixArray[26] = 12'h000;
iconPixArray[27] = 12'h000;
iconPixArray[28] = 12'h000;
iconPixArray[29] = 12'h000;
iconPixArray[30] = 12'h000;
iconPixArray[31] = 12'h000;
iconPixArray[32] = 12'h000;
iconPixArray[33] = 12'h000;
iconPixArray[34] = 12'h000;
iconPixArray[35] = 12'h000;
iconPixArray[36] = 12'h000;
iconPixArray[37] = 12'h000;
iconPixArray[38] = 12'h000;
iconPixArray[39] = 12'h000;
iconPixArray[40] = 12'h000;
iconPixArray[41] = 12'h000;
iconPixArray[42] = 12'h000;
iconPixArray[43] = 12'h000;
iconPixArray[44] = 12'h000;
iconPixArray[45] = 12'h000;
iconPixArray[46] = 12'h000;
iconPixArray[47] = 12'h000;
iconPixArray[48] = 12'h000;
iconPixArray[49] = 12'h000;
iconPixArray[50] = 12'h000;
iconPixArray[51] = 12'h000;
iconPixArray[52] = 12'h000;
iconPixArray[53] = 12'h000;
iconPixArray[54] = 12'h000;
iconPixArray[55] = 12'h000;
iconPixArray[56] = 12'h000;
iconPixArray[57] = 12'h000;
iconPixArray[58] = 12'h000;
iconPixArray[59] = 12'h000;
iconPixArray[60] = 12'h000;
iconPixArray[61] = 12'h000;
iconPixArray[62] = 12'h000;
iconPixArray[63] = 12'h000;
iconPixArray[64] = 12'h000;
iconPixArray[65] = 12'h000;
iconPixArray[66] = 12'h000;
iconPixArray[67] = 12'h000;
iconPixArray[68] = 12'h000;
iconPixArray[69] = 12'h000;
iconPixArray[70] = 12'h000;
iconPixArray[71] = 12'h000;
iconPixArray[72] = 12'h000;
iconPixArray[73] = 12'h000;
iconPixArray[74] = 12'h000;
iconPixArray[75] = 12'h000;
iconPixArray[76] = 12'h000;
iconPixArray[77] = 12'h000;
iconPixArray[78] = 12'h000;
iconPixArray[79] = 12'h000;
iconPixArray[80] = 12'h000;
iconPixArray[81] = 12'h000;
iconPixArray[82] = 12'h000;
iconPixArray[83] = 12'h000;
iconPixArray[84] = 12'h000;
iconPixArray[85] = 12'h000;
iconPixArray[86] = 12'h000;
iconPixArray[87] = 12'h000;
iconPixArray[88] = 12'h000;
iconPixArray[89] = 12'h000;
iconPixArray[90] = 12'h000;
iconPixArray[91] = 12'h133;
iconPixArray[92] = 12'h112;
iconPixArray[93] = 12'h000;
iconPixArray[94] = 12'h001;
iconPixArray[95] = 12'h000;
iconPixArray[96] = 12'h000;
iconPixArray[97] = 12'h000;
iconPixArray[98] = 12'h000;
iconPixArray[99] = 12'h000;
iconPixArray[100] = 12'h000;
iconPixArray[101] = 12'h000;
iconPixArray[102] = 12'h000;
iconPixArray[103] = 12'h000;
iconPixArray[104] = 12'h000;
iconPixArray[105] = 12'h000;
iconPixArray[106] = 12'h000;
iconPixArray[107] = 12'h000;
iconPixArray[108] = 12'h000;
iconPixArray[109] = 12'h000;
iconPixArray[110] = 12'h000;
iconPixArray[111] = 12'h000;
iconPixArray[112] = 12'h000;
iconPixArray[113] = 12'h000;
iconPixArray[114] = 12'h000;
iconPixArray[115] = 12'h000;
iconPixArray[116] = 12'h000;
iconPixArray[117] = 12'h000;
iconPixArray[118] = 12'h000;
iconPixArray[119] = 12'h000;
iconPixArray[120] = 12'h123;
iconPixArray[121] = 12'h000;
iconPixArray[122] = 12'h358;
iconPixArray[123] = 12'h6B0;
iconPixArray[124] = 12'h8F6;
iconPixArray[125] = 12'h7E5;
iconPixArray[126] = 12'h001;
iconPixArray[127] = 12'h000;
iconPixArray[128] = 12'h000;
iconPixArray[129] = 12'h000;
iconPixArray[130] = 12'h000;
iconPixArray[131] = 12'h000;
iconPixArray[132] = 12'h000;
iconPixArray[133] = 12'h000;
iconPixArray[134] = 12'h000;
iconPixArray[135] = 12'h000;
iconPixArray[136] = 12'h000;
iconPixArray[137] = 12'h000;
iconPixArray[138] = 12'h000;
iconPixArray[139] = 12'h000;
iconPixArray[140] = 12'h000;
iconPixArray[141] = 12'h000;
iconPixArray[142] = 12'h000;
iconPixArray[143] = 12'h000;
iconPixArray[144] = 12'h000;
iconPixArray[145] = 12'h000;
iconPixArray[146] = 12'h000;
iconPixArray[147] = 12'h000;
iconPixArray[148] = 12'h000;
iconPixArray[149] = 12'h001;
iconPixArray[150] = 12'h000;
iconPixArray[151] = 12'h358;
iconPixArray[152] = 12'h111;
iconPixArray[153] = 12'hD96;
iconPixArray[154] = 12'h469;
iconPixArray[155] = 12'h6AF;
iconPixArray[156] = 12'h6AF;
iconPixArray[157] = 12'h358;
iconPixArray[158] = 12'h123;
iconPixArray[159] = 12'h000;
iconPixArray[160] = 12'h000;
iconPixArray[161] = 12'h000;
iconPixArray[162] = 12'h000;
iconPixArray[163] = 12'h000;
iconPixArray[164] = 12'h000;
iconPixArray[165] = 12'h000;
iconPixArray[166] = 12'h000;
iconPixArray[167] = 12'h000;
iconPixArray[168] = 12'h000;
iconPixArray[169] = 12'h000;
iconPixArray[170] = 12'h000;
iconPixArray[171] = 12'h000;
iconPixArray[172] = 12'h000;
iconPixArray[173] = 12'h000;
iconPixArray[174] = 12'h000;
iconPixArray[175] = 12'h000;
iconPixArray[176] = 12'h000;
iconPixArray[177] = 12'h000;
iconPixArray[178] = 12'h000;
iconPixArray[179] = 12'h000;
iconPixArray[180] = 12'h011;
iconPixArray[181] = 12'h48C;
iconPixArray[182] = 12'hD84;
iconPixArray[183] = 12'h0FE;
iconPixArray[184] = 12'h6AF;
iconPixArray[185] = 12'h6AF;
iconPixArray[186] = 12'h6AF;
iconPixArray[187] = 12'h6AF;
iconPixArray[188] = 12'h6AF;
iconPixArray[189] = 12'h47A;
iconPixArray[190] = 12'h011;
iconPixArray[191] = 12'h000;
iconPixArray[192] = 12'h000;
iconPixArray[193] = 12'h000;
iconPixArray[194] = 12'h000;
iconPixArray[195] = 12'h000;
iconPixArray[196] = 12'h000;
iconPixArray[197] = 12'h000;
iconPixArray[198] = 12'h000;
iconPixArray[199] = 12'h000;
iconPixArray[200] = 12'h000;
iconPixArray[201] = 12'h000;
iconPixArray[202] = 12'h000;
iconPixArray[203] = 12'h000;
iconPixArray[204] = 12'h000;
iconPixArray[205] = 12'h000;
iconPixArray[206] = 12'h000;
iconPixArray[207] = 12'h000;
iconPixArray[208] = 12'h000;
iconPixArray[209] = 12'h000;
iconPixArray[210] = 12'h111;
iconPixArray[211] = 12'h000;
iconPixArray[212] = 12'hEB8;
iconPixArray[213] = 12'h0DC;
iconPixArray[214] = 12'h6AF;
iconPixArray[215] = 12'h6AF;
iconPixArray[216] = 12'h6AF;
iconPixArray[217] = 12'h6AF;
iconPixArray[218] = 12'h6AF;
iconPixArray[219] = 12'h6AF;
iconPixArray[220] = 12'h57B;
iconPixArray[221] = 12'h36A;
iconPixArray[222] = 12'h000;
iconPixArray[223] = 12'h000;
iconPixArray[224] = 12'h000;
iconPixArray[225] = 12'h000;
iconPixArray[226] = 12'h000;
iconPixArray[227] = 12'h000;
iconPixArray[228] = 12'h000;
iconPixArray[229] = 12'h000;
iconPixArray[230] = 12'h000;
iconPixArray[231] = 12'h000;
iconPixArray[232] = 12'h000;
iconPixArray[233] = 12'h000;
iconPixArray[234] = 12'h000;
iconPixArray[235] = 12'h000;
iconPixArray[236] = 12'h000;
iconPixArray[237] = 12'h000;
iconPixArray[238] = 12'h000;
iconPixArray[239] = 12'h000;
iconPixArray[240] = 12'h000;
iconPixArray[241] = 12'h125;
iconPixArray[242] = 12'h245;
iconPixArray[243] = 12'h6AF;
iconPixArray[244] = 12'h6AF;
iconPixArray[245] = 12'h6AF;
iconPixArray[246] = 12'h6AF;
iconPixArray[247] = 12'h6AF;
iconPixArray[248] = 12'h6AF;
iconPixArray[249] = 12'h6AF;
iconPixArray[250] = 12'h6AF;
iconPixArray[251] = 12'h6AF;
iconPixArray[252] = 12'h111;
iconPixArray[253] = 12'h000;
iconPixArray[254] = 12'h000;
iconPixArray[255] = 12'h000;
iconPixArray[256] = 12'h000;
iconPixArray[257] = 12'h000;
iconPixArray[258] = 12'h000;
iconPixArray[259] = 12'h000;
iconPixArray[260] = 12'h000;
iconPixArray[261] = 12'h000;
iconPixArray[262] = 12'h000;
iconPixArray[263] = 12'h000;
iconPixArray[264] = 12'h000;
iconPixArray[265] = 12'h000;
iconPixArray[266] = 12'h000;
iconPixArray[267] = 12'h000;
iconPixArray[268] = 12'h000;
iconPixArray[269] = 12'h000;
iconPixArray[270] = 12'h000;
iconPixArray[271] = 12'h000;
iconPixArray[272] = 12'h123;
iconPixArray[273] = 12'h6D3;
iconPixArray[274] = 12'h234;
iconPixArray[275] = 12'h212;
iconPixArray[276] = 12'hC97;
iconPixArray[277] = 12'hF37;
iconPixArray[278] = 12'hD14;
iconPixArray[279] = 12'h38D;
iconPixArray[280] = 12'hB4E;
iconPixArray[281] = 12'h6AF;
iconPixArray[282] = 12'h6AF;
iconPixArray[283] = 12'h6AF;
iconPixArray[284] = 12'h6C2;
iconPixArray[285] = 12'h011;
iconPixArray[286] = 12'h000;
iconPixArray[287] = 12'h000;
iconPixArray[288] = 12'h000;
iconPixArray[289] = 12'h000;
iconPixArray[290] = 12'h000;
iconPixArray[291] = 12'h000;
iconPixArray[292] = 12'h000;
iconPixArray[293] = 12'h000;
iconPixArray[294] = 12'h000;
iconPixArray[295] = 12'h000;
iconPixArray[296] = 12'h000;
iconPixArray[297] = 12'h000;
iconPixArray[298] = 12'h000;
iconPixArray[299] = 12'h000;
iconPixArray[300] = 12'h000;
iconPixArray[301] = 12'h000;
iconPixArray[302] = 12'h000;
iconPixArray[303] = 12'h123;
iconPixArray[304] = 12'hC84;
iconPixArray[305] = 12'hB5F;
iconPixArray[306] = 12'h69E;
iconPixArray[307] = 12'h136;
iconPixArray[308] = 12'hF14;
iconPixArray[309] = 12'h777;
iconPixArray[310] = 12'hFFF;
iconPixArray[311] = 12'h778;
iconPixArray[312] = 12'h709;
iconPixArray[313] = 12'h223;
iconPixArray[314] = 12'h6AF;
iconPixArray[315] = 12'h458;
iconPixArray[316] = 12'h6C1;
iconPixArray[317] = 12'h001;
iconPixArray[318] = 12'h000;
iconPixArray[319] = 12'h000;
iconPixArray[320] = 12'h000;
iconPixArray[321] = 12'h000;
iconPixArray[322] = 12'h000;
iconPixArray[323] = 12'h000;
iconPixArray[324] = 12'h000;
iconPixArray[325] = 12'h000;
iconPixArray[326] = 12'h000;
iconPixArray[327] = 12'h000;
iconPixArray[328] = 12'h000;
iconPixArray[329] = 12'h000;
iconPixArray[330] = 12'h000;
iconPixArray[331] = 12'h000;
iconPixArray[332] = 12'h000;
iconPixArray[333] = 12'h000;
iconPixArray[334] = 12'h123;
iconPixArray[335] = 12'h91A;
iconPixArray[336] = 12'hC72;
iconPixArray[337] = 12'h6AF;
iconPixArray[338] = 12'h357;
iconPixArray[339] = 12'h9E4;
iconPixArray[340] = 12'hFFF;
iconPixArray[341] = 12'hFFF;
iconPixArray[342] = 12'hFFF;
iconPixArray[343] = 12'hFFF;
iconPixArray[344] = 12'hC03;
iconPixArray[345] = 12'h58C;
iconPixArray[346] = 12'h6AF;
iconPixArray[347] = 12'h58C;
iconPixArray[348] = 12'h000;
iconPixArray[349] = 12'h000;
iconPixArray[350] = 12'h000;
iconPixArray[351] = 12'h000;
iconPixArray[352] = 12'h000;
iconPixArray[353] = 12'h000;
iconPixArray[354] = 12'h000;
iconPixArray[355] = 12'h000;
iconPixArray[356] = 12'h000;
iconPixArray[357] = 12'h000;
iconPixArray[358] = 12'h000;
iconPixArray[359] = 12'h000;
iconPixArray[360] = 12'h000;
iconPixArray[361] = 12'h000;
iconPixArray[362] = 12'h000;
iconPixArray[363] = 12'h000;
iconPixArray[364] = 12'h000;
iconPixArray[365] = 12'h123;
iconPixArray[366] = 12'h6C1;
iconPixArray[367] = 12'h9F7;
iconPixArray[368] = 12'h6AF;
iconPixArray[369] = 12'h6AF;
iconPixArray[370] = 12'h8F7;
iconPixArray[371] = 12'h8C0;
iconPixArray[372] = 12'hFFF;
iconPixArray[373] = 12'hFFF;
iconPixArray[374] = 12'hFFF;
iconPixArray[375] = 12'hFFF;
iconPixArray[376] = 12'hCCC;
iconPixArray[377] = 12'hF4B;
iconPixArray[378] = 12'h469;
iconPixArray[379] = 12'hA3D;
iconPixArray[380] = 12'h113;
iconPixArray[381] = 12'h000;
iconPixArray[382] = 12'h000;
iconPixArray[383] = 12'h000;
iconPixArray[384] = 12'h000;
iconPixArray[385] = 12'h000;
iconPixArray[386] = 12'h000;
iconPixArray[387] = 12'h000;
iconPixArray[388] = 12'h000;
iconPixArray[389] = 12'h000;
iconPixArray[390] = 12'h000;
iconPixArray[391] = 12'h000;
iconPixArray[392] = 12'h100;
iconPixArray[393] = 12'h500;
iconPixArray[394] = 12'h500;
iconPixArray[395] = 12'h100;
iconPixArray[396] = 12'h001;
iconPixArray[397] = 12'h235;
iconPixArray[398] = 12'h358;
iconPixArray[399] = 12'h6AF;
iconPixArray[400] = 12'h6AF;
iconPixArray[401] = 12'h6AF;
iconPixArray[402] = 12'h9F7;
iconPixArray[403] = 12'h49E;
iconPixArray[404] = 12'hBBB;
iconPixArray[405] = 12'hFFF;
iconPixArray[406] = 12'hFFF;
iconPixArray[407] = 12'hFFF;
iconPixArray[408] = 12'hC16;
iconPixArray[409] = 12'hA2B;
iconPixArray[410] = 12'hC73;
iconPixArray[411] = 12'h000;
iconPixArray[412] = 12'h000;
iconPixArray[413] = 12'h000;
iconPixArray[414] = 12'h000;
iconPixArray[415] = 12'h000;
iconPixArray[416] = 12'h000;
iconPixArray[417] = 12'h000;
iconPixArray[418] = 12'h000;
iconPixArray[419] = 12'h000;
iconPixArray[420] = 12'h000;
iconPixArray[421] = 12'h000;
iconPixArray[422] = 12'h200;
iconPixArray[423] = 12'h000;
iconPixArray[424] = 12'hC00;
iconPixArray[425] = 12'h200;
iconPixArray[426] = 12'h200;
iconPixArray[427] = 12'hE00;
iconPixArray[428] = 12'h000;
iconPixArray[429] = 12'h112;
iconPixArray[430] = 12'h57B;
iconPixArray[431] = 12'h7BF;
iconPixArray[432] = 12'h0EB;
iconPixArray[433] = 12'h28F;
iconPixArray[434] = 12'hB4E;
iconPixArray[435] = 12'hF02;
iconPixArray[436] = 12'hC15;
iconPixArray[437] = 12'hEEE;
iconPixArray[438] = 12'h000;
iconPixArray[439] = 12'h48C;
iconPixArray[440] = 12'hF01;
iconPixArray[441] = 12'h5AE;
iconPixArray[442] = 12'h235;
iconPixArray[443] = 12'h000;
iconPixArray[444] = 12'h000;
iconPixArray[445] = 12'h000;
iconPixArray[446] = 12'h000;
iconPixArray[447] = 12'h000;
iconPixArray[448] = 12'h000;
iconPixArray[449] = 12'h000;
iconPixArray[450] = 12'h000;
iconPixArray[451] = 12'h000;
iconPixArray[452] = 12'h000;
iconPixArray[453] = 12'h000;
iconPixArray[454] = 12'h000;
iconPixArray[455] = 12'hB00;
iconPixArray[456] = 12'hF00;
iconPixArray[457] = 12'hF00;
iconPixArray[458] = 12'h700;
iconPixArray[459] = 12'h900;
iconPixArray[460] = 12'hB4D;
iconPixArray[461] = 12'h346;
iconPixArray[462] = 12'hB86;
iconPixArray[463] = 12'h148;
iconPixArray[464] = 12'h555;
iconPixArray[465] = 12'hFF0;
iconPixArray[466] = 12'h8D2;
iconPixArray[467] = 12'h0ED;
iconPixArray[468] = 12'hB18;
iconPixArray[469] = 12'h7AD;
iconPixArray[470] = 12'h333;
iconPixArray[471] = 12'h520;
iconPixArray[472] = 12'hDA6;
iconPixArray[473] = 12'hA3D;
iconPixArray[474] = 12'h123;
iconPixArray[475] = 12'h000;
iconPixArray[476] = 12'h000;
iconPixArray[477] = 12'h000;
iconPixArray[478] = 12'h000;
iconPixArray[479] = 12'h000;
iconPixArray[480] = 12'h000;
iconPixArray[481] = 12'h000;
iconPixArray[482] = 12'h000;
iconPixArray[483] = 12'h000;
iconPixArray[484] = 12'h000;
iconPixArray[485] = 12'h100;
iconPixArray[486] = 12'hA00;
iconPixArray[487] = 12'hF00;
iconPixArray[488] = 12'hF00;
iconPixArray[489] = 12'h800;
iconPixArray[490] = 12'hD00;
iconPixArray[491] = 12'h434;
iconPixArray[492] = 12'hC61;
iconPixArray[493] = 12'h3FA;
iconPixArray[494] = 12'hAE1;
iconPixArray[495] = 12'hFFF;
iconPixArray[496] = 12'hFFF;
iconPixArray[497] = 12'hFFF;
iconPixArray[498] = 12'h777;
iconPixArray[499] = 12'h7F7;
iconPixArray[500] = 12'h69E;
iconPixArray[501] = 12'h6AF;
iconPixArray[502] = 12'h6AF;
iconPixArray[503] = 12'h47A;
iconPixArray[504] = 12'h59E;
iconPixArray[505] = 12'h122;
iconPixArray[506] = 12'h000;
iconPixArray[507] = 12'h000;
iconPixArray[508] = 12'h000;
iconPixArray[509] = 12'h000;
iconPixArray[510] = 12'h000;
iconPixArray[511] = 12'h000;
iconPixArray[512] = 12'h000;
iconPixArray[513] = 12'h000;
iconPixArray[514] = 12'h000;
iconPixArray[515] = 12'h000;
iconPixArray[516] = 12'h400;
iconPixArray[517] = 12'h900;
iconPixArray[518] = 12'h100;
iconPixArray[519] = 12'hF00;
iconPixArray[520] = 12'hF00;
iconPixArray[521] = 12'hE00;
iconPixArray[522] = 12'h000;
iconPixArray[523] = 12'h58C;
iconPixArray[524] = 12'h6AF;
iconPixArray[525] = 12'h68B;
iconPixArray[526] = 12'hCCC;
iconPixArray[527] = 12'hFFF;
iconPixArray[528] = 12'hFFF;
iconPixArray[529] = 12'hFFF;
iconPixArray[530] = 12'hFFF;
iconPixArray[531] = 12'hD39;
iconPixArray[532] = 12'hB4E;
iconPixArray[533] = 12'h6AF;
iconPixArray[534] = 12'h59D;
iconPixArray[535] = 12'h0FE;
iconPixArray[536] = 12'h000;
iconPixArray[537] = 12'h000;
iconPixArray[538] = 12'h000;
iconPixArray[539] = 12'h000;
iconPixArray[540] = 12'h000;
iconPixArray[541] = 12'h000;
iconPixArray[542] = 12'h000;
iconPixArray[543] = 12'h000;
iconPixArray[544] = 12'h000;
iconPixArray[545] = 12'h000;
iconPixArray[546] = 12'h000;
iconPixArray[547] = 12'h000;
iconPixArray[548] = 12'h000;
iconPixArray[549] = 12'h600;
iconPixArray[550] = 12'hF00;
iconPixArray[551] = 12'hF00;
iconPixArray[552] = 12'h300;
iconPixArray[553] = 12'h100;
iconPixArray[554] = 12'h8F7;
iconPixArray[555] = 12'h6AF;
iconPixArray[556] = 12'h6AF;
iconPixArray[557] = 12'hC61;
iconPixArray[558] = 12'h333;
iconPixArray[559] = 12'hFFF;
iconPixArray[560] = 12'hFFF;
iconPixArray[561] = 12'hFFF;
iconPixArray[562] = 12'hDDD;
iconPixArray[563] = 12'h8D1;
iconPixArray[564] = 12'h212;
iconPixArray[565] = 12'h58C;
iconPixArray[566] = 12'hFEC;
iconPixArray[567] = 12'h000;
iconPixArray[568] = 12'h000;
iconPixArray[569] = 12'h000;
iconPixArray[570] = 12'h000;
iconPixArray[571] = 12'h000;
iconPixArray[572] = 12'h000;
iconPixArray[573] = 12'h000;
iconPixArray[574] = 12'h000;
iconPixArray[575] = 12'h000;
iconPixArray[576] = 12'h000;
iconPixArray[577] = 12'h000;
iconPixArray[578] = 12'h000;
iconPixArray[579] = 12'h200;
iconPixArray[580] = 12'h600;
iconPixArray[581] = 12'hD00;
iconPixArray[582] = 12'hF00;
iconPixArray[583] = 12'h000;
iconPixArray[584] = 12'hD00;
iconPixArray[585] = 12'h8C2;
iconPixArray[586] = 12'h458;
iconPixArray[587] = 12'h6AF;
iconPixArray[588] = 12'h6AF;
iconPixArray[589] = 12'h358;
iconPixArray[590] = 12'h38D;
iconPixArray[591] = 12'h000;
iconPixArray[592] = 12'hFFF;
iconPixArray[593] = 12'hEEE;
iconPixArray[594] = 12'hABD;
iconPixArray[595] = 12'h83D;
iconPixArray[596] = 12'h57B;
iconPixArray[597] = 12'hECA;
iconPixArray[598] = 12'h000;
iconPixArray[599] = 12'h000;
iconPixArray[600] = 12'h000;
iconPixArray[601] = 12'h000;
iconPixArray[602] = 12'h000;
iconPixArray[603] = 12'h000;
iconPixArray[604] = 12'h000;
iconPixArray[605] = 12'h000;
iconPixArray[606] = 12'h000;
iconPixArray[607] = 12'h000;
iconPixArray[608] = 12'h000;
iconPixArray[609] = 12'h000;
iconPixArray[610] = 12'h000;
iconPixArray[611] = 12'h000;
iconPixArray[612] = 12'h700;
iconPixArray[613] = 12'hF00;
iconPixArray[614] = 12'hE00;
iconPixArray[615] = 12'hE00;
iconPixArray[616] = 12'h211;
iconPixArray[617] = 12'h469;
iconPixArray[618] = 12'h6AF;
iconPixArray[619] = 12'h6AF;
iconPixArray[620] = 12'h6AF;
iconPixArray[621] = 12'h6AF;
iconPixArray[622] = 12'hC3B;
iconPixArray[623] = 12'h4A0;
iconPixArray[624] = 12'hD3A;
iconPixArray[625] = 12'hC17;
iconPixArray[626] = 12'h82D;
iconPixArray[627] = 12'hC50;
iconPixArray[628] = 12'h00F;
iconPixArray[629] = 12'h000;
iconPixArray[630] = 12'h000;
iconPixArray[631] = 12'h000;
iconPixArray[632] = 12'h000;
iconPixArray[633] = 12'h000;
iconPixArray[634] = 12'h000;
iconPixArray[635] = 12'h000;
iconPixArray[636] = 12'h000;
iconPixArray[637] = 12'h000;
iconPixArray[638] = 12'h000;
iconPixArray[639] = 12'h000;
iconPixArray[640] = 12'h000;
iconPixArray[641] = 12'h000;
iconPixArray[642] = 12'h000;
iconPixArray[643] = 12'h200;
iconPixArray[644] = 12'h400;
iconPixArray[645] = 12'h800;
iconPixArray[646] = 12'h100;
iconPixArray[647] = 12'h000;
iconPixArray[648] = 12'h7D4;
iconPixArray[649] = 12'h6AF;
iconPixArray[650] = 12'h6AF;
iconPixArray[651] = 12'h6AF;
iconPixArray[652] = 12'h6AF;
iconPixArray[653] = 12'h6AF;
iconPixArray[654] = 12'h6AF;
iconPixArray[655] = 12'h69E;
iconPixArray[656] = 12'hD73;
iconPixArray[657] = 12'h346;
iconPixArray[658] = 12'h69D;
iconPixArray[659] = 12'h58B;
iconPixArray[660] = 12'h000;
iconPixArray[661] = 12'h000;
iconPixArray[662] = 12'h000;
iconPixArray[663] = 12'h000;
iconPixArray[664] = 12'h000;
iconPixArray[665] = 12'h000;
iconPixArray[666] = 12'h000;
iconPixArray[667] = 12'h000;
iconPixArray[668] = 12'h000;
iconPixArray[669] = 12'h000;
iconPixArray[670] = 12'h000;
iconPixArray[671] = 12'h000;
iconPixArray[672] = 12'h000;
iconPixArray[673] = 12'h000;
iconPixArray[674] = 12'h300;
iconPixArray[675] = 12'h000;
iconPixArray[676] = 12'h000;
iconPixArray[677] = 12'h200;
iconPixArray[678] = 12'h000;
iconPixArray[679] = 12'h001;
iconPixArray[680] = 12'h8F7;
iconPixArray[681] = 12'h346;
iconPixArray[682] = 12'h6AF;
iconPixArray[683] = 12'h6AF;
iconPixArray[684] = 12'h6AF;
iconPixArray[685] = 12'h6AF;
iconPixArray[686] = 12'h6AF;
iconPixArray[687] = 12'h6AF;
iconPixArray[688] = 12'h6AF;
iconPixArray[689] = 12'h369;
iconPixArray[690] = 12'h512;
iconPixArray[691] = 12'h500;
iconPixArray[692] = 12'h500;
iconPixArray[693] = 12'h000;
iconPixArray[694] = 12'h000;
iconPixArray[695] = 12'h000;
iconPixArray[696] = 12'h000;
iconPixArray[697] = 12'h000;
iconPixArray[698] = 12'h000;
iconPixArray[699] = 12'h000;
iconPixArray[700] = 12'h000;
iconPixArray[701] = 12'h000;
iconPixArray[702] = 12'h000;
iconPixArray[703] = 12'h000;
iconPixArray[704] = 12'h000;
iconPixArray[705] = 12'h000;
iconPixArray[706] = 12'h000;
iconPixArray[707] = 12'h000;
iconPixArray[708] = 12'h000;
iconPixArray[709] = 12'h000;
iconPixArray[710] = 12'h000;
iconPixArray[711] = 12'h000;
iconPixArray[712] = 12'h011;
iconPixArray[713] = 12'h6B2;
iconPixArray[714] = 12'h335;
iconPixArray[715] = 12'h6AF;
iconPixArray[716] = 12'h6AF;
iconPixArray[717] = 12'h6AF;
iconPixArray[718] = 12'h6AF;
iconPixArray[719] = 12'h6AF;
iconPixArray[720] = 12'hD96;
iconPixArray[721] = 12'h200;
iconPixArray[722] = 12'hB00;
iconPixArray[723] = 12'h800;
iconPixArray[724] = 12'h800;
iconPixArray[725] = 12'h000;
iconPixArray[726] = 12'h000;
iconPixArray[727] = 12'h000;
iconPixArray[728] = 12'h000;
iconPixArray[729] = 12'h000;
iconPixArray[730] = 12'h000;
iconPixArray[731] = 12'h000;
iconPixArray[732] = 12'h000;
iconPixArray[733] = 12'h000;
iconPixArray[734] = 12'h000;
iconPixArray[735] = 12'h000;
iconPixArray[736] = 12'h000;
iconPixArray[737] = 12'h000;
iconPixArray[738] = 12'h000;
iconPixArray[739] = 12'h000;
iconPixArray[740] = 12'h000;
iconPixArray[741] = 12'h000;
iconPixArray[742] = 12'h000;
iconPixArray[743] = 12'h000;
iconPixArray[744] = 12'h000;
iconPixArray[745] = 12'h112;
iconPixArray[746] = 12'h112;
iconPixArray[747] = 12'h0ED;
iconPixArray[748] = 12'h6AF;
iconPixArray[749] = 12'h6AF;
iconPixArray[750] = 12'hEB8;
iconPixArray[751] = 12'hA3C;
iconPixArray[752] = 12'h000;
iconPixArray[753] = 12'h600;
iconPixArray[754] = 12'hB00;
iconPixArray[755] = 12'hF00;
iconPixArray[756] = 12'hE00;
iconPixArray[757] = 12'h000;
iconPixArray[758] = 12'h000;
iconPixArray[759] = 12'h000;
iconPixArray[760] = 12'h000;
iconPixArray[761] = 12'h000;
iconPixArray[762] = 12'h000;
iconPixArray[763] = 12'h000;
iconPixArray[764] = 12'h000;
iconPixArray[765] = 12'h000;
iconPixArray[766] = 12'h000;
iconPixArray[767] = 12'h000;
iconPixArray[768] = 12'h000;
iconPixArray[769] = 12'h000;
iconPixArray[770] = 12'h000;
iconPixArray[771] = 12'h000;
iconPixArray[772] = 12'h000;
iconPixArray[773] = 12'h000;
iconPixArray[774] = 12'h000;
iconPixArray[775] = 12'h000;
iconPixArray[776] = 12'h000;
iconPixArray[777] = 12'h000;
iconPixArray[778] = 12'h112;
iconPixArray[779] = 12'h000;
iconPixArray[780] = 12'h0DC;
iconPixArray[781] = 12'hEA7;
iconPixArray[782] = 12'h546;
iconPixArray[783] = 12'h100;
iconPixArray[784] = 12'hF00;
iconPixArray[785] = 12'hD00;
iconPixArray[786] = 12'hF00;
iconPixArray[787] = 12'hD00;
iconPixArray[788] = 12'h200;
iconPixArray[789] = 12'h000;
iconPixArray[790] = 12'h000;
iconPixArray[791] = 12'h000;
iconPixArray[792] = 12'h000;
iconPixArray[793] = 12'h000;
iconPixArray[794] = 12'h000;
iconPixArray[795] = 12'h000;
iconPixArray[796] = 12'h000;
iconPixArray[797] = 12'h000;
iconPixArray[798] = 12'h000;
iconPixArray[799] = 12'h000;
iconPixArray[800] = 12'h000;
iconPixArray[801] = 12'h000;
iconPixArray[802] = 12'h000;
iconPixArray[803] = 12'h000;
iconPixArray[804] = 12'h000;
iconPixArray[805] = 12'h000;
iconPixArray[806] = 12'h000;
iconPixArray[807] = 12'h000;
iconPixArray[808] = 12'h000;
iconPixArray[809] = 12'h000;
iconPixArray[810] = 12'h000;
iconPixArray[811] = 12'h112;
iconPixArray[812] = 12'hEB9;
iconPixArray[813] = 12'h311;
iconPixArray[814] = 12'h100;
iconPixArray[815] = 12'h800;
iconPixArray[816] = 12'hF00;
iconPixArray[817] = 12'hF00;
iconPixArray[818] = 12'hF00;
iconPixArray[819] = 12'h000;
iconPixArray[820] = 12'h000;
iconPixArray[821] = 12'h000;
iconPixArray[822] = 12'h000;
iconPixArray[823] = 12'h000;
iconPixArray[824] = 12'h000;
iconPixArray[825] = 12'h000;
iconPixArray[826] = 12'h000;
iconPixArray[827] = 12'h000;
iconPixArray[828] = 12'h000;
iconPixArray[829] = 12'h000;
iconPixArray[830] = 12'h000;
iconPixArray[831] = 12'h000;
iconPixArray[832] = 12'h000;
iconPixArray[833] = 12'h000;
iconPixArray[834] = 12'h000;
iconPixArray[835] = 12'h000;
iconPixArray[836] = 12'h000;
iconPixArray[837] = 12'h000;
iconPixArray[838] = 12'h000;
iconPixArray[839] = 12'h000;
iconPixArray[840] = 12'h000;
iconPixArray[841] = 12'h000;
iconPixArray[842] = 12'h000;
iconPixArray[843] = 12'h000;
iconPixArray[844] = 12'h111;
iconPixArray[845] = 12'h000;
iconPixArray[846] = 12'hE00;
iconPixArray[847] = 12'hF00;
iconPixArray[848] = 12'hF00;
iconPixArray[849] = 12'hE00;
iconPixArray[850] = 12'h000;
iconPixArray[851] = 12'h200;
iconPixArray[852] = 12'h100;
iconPixArray[853] = 12'h000;
iconPixArray[854] = 12'h000;
iconPixArray[855] = 12'h000;
iconPixArray[856] = 12'h000;
iconPixArray[857] = 12'h000;
iconPixArray[858] = 12'h000;
iconPixArray[859] = 12'h000;
iconPixArray[860] = 12'h000;
iconPixArray[861] = 12'h000;
iconPixArray[862] = 12'h000;
iconPixArray[863] = 12'h000;
iconPixArray[864] = 12'h000;
iconPixArray[865] = 12'h000;
iconPixArray[866] = 12'h000;
iconPixArray[867] = 12'h000;
iconPixArray[868] = 12'h000;
iconPixArray[869] = 12'h000;
iconPixArray[870] = 12'h000;
iconPixArray[871] = 12'h000;
iconPixArray[872] = 12'h000;
iconPixArray[873] = 12'h000;
iconPixArray[874] = 12'h000;
iconPixArray[875] = 12'h000;
iconPixArray[876] = 12'h100;
iconPixArray[877] = 12'h100;
iconPixArray[878] = 12'hF00;
iconPixArray[879] = 12'hF00;
iconPixArray[880] = 12'hC00;
iconPixArray[881] = 12'h000;
iconPixArray[882] = 12'h000;
iconPixArray[883] = 12'h300;
iconPixArray[884] = 12'h000;
iconPixArray[885] = 12'h000;
iconPixArray[886] = 12'h000;
iconPixArray[887] = 12'h000;
iconPixArray[888] = 12'h000;
iconPixArray[889] = 12'h000;
iconPixArray[890] = 12'h000;
iconPixArray[891] = 12'h000;
iconPixArray[892] = 12'h000;
iconPixArray[893] = 12'h000;
iconPixArray[894] = 12'h000;
iconPixArray[895] = 12'h000;
iconPixArray[896] = 12'h000;
iconPixArray[897] = 12'h000;
iconPixArray[898] = 12'h000;
iconPixArray[899] = 12'h000;
iconPixArray[900] = 12'h000;
iconPixArray[901] = 12'h000;
iconPixArray[902] = 12'h000;
iconPixArray[903] = 12'h000;
iconPixArray[904] = 12'h000;
iconPixArray[905] = 12'h000;
iconPixArray[906] = 12'h000;
iconPixArray[907] = 12'h000;
iconPixArray[908] = 12'h100;
iconPixArray[909] = 12'h700;
iconPixArray[910] = 12'h700;
iconPixArray[911] = 12'h500;
iconPixArray[912] = 12'h200;
iconPixArray[913] = 12'h300;
iconPixArray[914] = 12'h000;
iconPixArray[915] = 12'h000;
iconPixArray[916] = 12'h000;
iconPixArray[917] = 12'h000;
iconPixArray[918] = 12'h000;
iconPixArray[919] = 12'h000;
iconPixArray[920] = 12'h000;
iconPixArray[921] = 12'h000;
iconPixArray[922] = 12'h000;
iconPixArray[923] = 12'h000;
iconPixArray[924] = 12'h000;
iconPixArray[925] = 12'h000;
iconPixArray[926] = 12'h000;
iconPixArray[927] = 12'h000;
iconPixArray[928] = 12'h000;
iconPixArray[929] = 12'h000;
iconPixArray[930] = 12'h000;
iconPixArray[931] = 12'h000;
iconPixArray[932] = 12'h000;
iconPixArray[933] = 12'h000;
iconPixArray[934] = 12'h000;
iconPixArray[935] = 12'h000;
iconPixArray[936] = 12'h000;
iconPixArray[937] = 12'h000;
iconPixArray[938] = 12'h000;
iconPixArray[939] = 12'h000;
iconPixArray[940] = 12'h000;
iconPixArray[941] = 12'hD00;
iconPixArray[942] = 12'h400;
iconPixArray[943] = 12'h200;
iconPixArray[944] = 12'h000;
iconPixArray[945] = 12'h000;
iconPixArray[946] = 12'h000;
iconPixArray[947] = 12'h000;
iconPixArray[948] = 12'h000;
iconPixArray[949] = 12'h000;
iconPixArray[950] = 12'h000;
iconPixArray[951] = 12'h000;
iconPixArray[952] = 12'h000;
iconPixArray[953] = 12'h000;
iconPixArray[954] = 12'h000;
iconPixArray[955] = 12'h000;
iconPixArray[956] = 12'h000;
iconPixArray[957] = 12'h000;
iconPixArray[958] = 12'h000;
iconPixArray[959] = 12'h000;
iconPixArray[960] = 12'h000;
iconPixArray[961] = 12'h000;
iconPixArray[962] = 12'h000;
iconPixArray[963] = 12'h000;
iconPixArray[964] = 12'h000;
iconPixArray[965] = 12'h000;
iconPixArray[966] = 12'h000;
iconPixArray[967] = 12'h000;
iconPixArray[968] = 12'h000;
iconPixArray[969] = 12'h000;
iconPixArray[970] = 12'h000;
iconPixArray[971] = 12'h000;
iconPixArray[972] = 12'h000;
iconPixArray[973] = 12'h300;
iconPixArray[974] = 12'h000;
iconPixArray[975] = 12'h000;
iconPixArray[976] = 12'h000;
iconPixArray[977] = 12'h000;
iconPixArray[978] = 12'h000;
iconPixArray[979] = 12'h000;
iconPixArray[980] = 12'h000;
iconPixArray[981] = 12'h000;
iconPixArray[982] = 12'h000;
iconPixArray[983] = 12'h000;
iconPixArray[984] = 12'h000;
iconPixArray[985] = 12'h000;
iconPixArray[986] = 12'h000;
iconPixArray[987] = 12'h000;
iconPixArray[988] = 12'h000;
iconPixArray[989] = 12'h000;
iconPixArray[990] = 12'h000;
iconPixArray[991] = 12'h000;
iconPixArray[992] = 12'h000;
iconPixArray[993] = 12'h000;
iconPixArray[994] = 12'h000;
iconPixArray[995] = 12'h000;
iconPixArray[996] = 12'h000;
iconPixArray[997] = 12'h000;
iconPixArray[998] = 12'h000;
iconPixArray[999] = 12'h000;
iconPixArray[1000] = 12'h000;
iconPixArray[1001] = 12'h000;
iconPixArray[1002] = 12'h000;
iconPixArray[1003] = 12'h000;
iconPixArray[1004] = 12'h000;
iconPixArray[1005] = 12'h000;
iconPixArray[1006] = 12'h000;
iconPixArray[1007] = 12'h000;
iconPixArray[1008] = 12'h000;
iconPixArray[1009] = 12'h000;
iconPixArray[1010] = 12'h000;
iconPixArray[1011] = 12'h000;
iconPixArray[1012] = 12'h000;
iconPixArray[1013] = 12'h000;
iconPixArray[1014] = 12'h000;
iconPixArray[1015] = 12'h000;
iconPixArray[1016] = 12'h000;
iconPixArray[1017] = 12'h000;
iconPixArray[1018] = 12'h000;
iconPixArray[1019] = 12'h000;
iconPixArray[1020] = 12'h000;
iconPixArray[1021] = 12'h000;
iconPixArray[1022] = 12'h000;
iconPixArray[1023] = 12'h000;
*/
/**********************************************
*****  Template file for the image array
*****  Produced from favicon.ico
***********************************************/
iconPixArray[256] = 12'h 00;
iconPixArray[257] = 12'h 00;
iconPixArray[258] = 12'h 00;
iconPixArray[259] = 12'h 00;
iconPixArray[260] = 12'h 00;
iconPixArray[261] = 12'h 00;
iconPixArray[262] = 12'h 00;
iconPixArray[263] = 12'h 00;
iconPixArray[264] = 12'h 00;
iconPixArray[265] = 12'h 00;
iconPixArray[266] = 12'h 00;
iconPixArray[267] = 12'h 00;
iconPixArray[268] = 12'h 00;
iconPixArray[269] = 12'h 00;
iconPixArray[270] = 12'h 00;
iconPixArray[271] = 12'h 00;
iconPixArray[272] = 12'h 00;
iconPixArray[273] = 12'h 00;
iconPixArray[274] = 12'h 00;
iconPixArray[275] = 12'h 00;
iconPixArray[276] = 12'h 00;
iconPixArray[277] = 12'h 00;
iconPixArray[278] = 12'h 00;
iconPixArray[279] = 12'h 00;
iconPixArray[280] = 12'h 00;
iconPixArray[281] = 12'h 00;
iconPixArray[282] = 12'h 00;
iconPixArray[283] = 12'h 00;
iconPixArray[284] = 12'h 11;
iconPixArray[285] = 12'h 11;
iconPixArray[286] = 12'h 11;
iconPixArray[287] = 12'h 01;
iconPixArray[288] = 12'h 00;
iconPixArray[289] = 12'h 00;
iconPixArray[290] = 12'h 00;
iconPixArray[291] = 12'h 00;
iconPixArray[292] = 12'h 00;
iconPixArray[293] = 12'h 00;
iconPixArray[294] = 12'h 00;
iconPixArray[295] = 12'h 00;
iconPixArray[296] = 12'h 00;
iconPixArray[297] = 12'h 00;
iconPixArray[298] = 12'h 11;
iconPixArray[299] = 12'h124;
iconPixArray[300] = 12'h37A;
iconPixArray[301] = 12'h59E;
iconPixArray[302] = 12'h369;
iconPixArray[303] = 12'h 00;
iconPixArray[304] = 12'h 00;
iconPixArray[305] = 12'h 00;
iconPixArray[306] = 12'h 00;
iconPixArray[307] = 12'h 00;
iconPixArray[308] = 12'h 00;
iconPixArray[309] = 12'h 00;
iconPixArray[310] = 12'h 00;
iconPixArray[311] = 12'h 00;
iconPixArray[312] = 12'h 00;
iconPixArray[313] = 12'h 12;
iconPixArray[314] = 12'h47B;
iconPixArray[315] = 12'h5AF;
iconPixArray[316] = 12'h5AF;
iconPixArray[317] = 12'h5AF;
iconPixArray[318] = 12'h135;
iconPixArray[319] = 12'h 00;
iconPixArray[320] = 12'h 00;
iconPixArray[321] = 12'h 00;
iconPixArray[322] = 12'h 00;
iconPixArray[323] = 12'h 00;
iconPixArray[324] = 12'h 00;
iconPixArray[325] = 12'h 00;
iconPixArray[326] = 12'h 00;
iconPixArray[327] = 12'h 01;
iconPixArray[328] = 12'h123;
iconPixArray[329] = 12'h47B;
iconPixArray[330] = 12'h567;
iconPixArray[331] = 12'h677;
iconPixArray[332] = 12'h47B;
iconPixArray[333] = 12'h59E;
iconPixArray[334] = 12'h 11;
iconPixArray[335] = 12'h 00;
iconPixArray[336] = 12'h 00;
iconPixArray[337] = 12'h 00;
iconPixArray[338] = 12'h 00;
iconPixArray[339] = 12'h 00;
iconPixArray[340] = 12'h 00;
iconPixArray[341] = 12'h 00;
iconPixArray[342] = 12'h 01;
iconPixArray[343] = 12'h123;
iconPixArray[344] = 12'h49E;
iconPixArray[345] = 12'h468;
iconPixArray[346] = 12'hFFF;
iconPixArray[347] = 12'hFFF;
iconPixArray[348] = 12'h568;
iconPixArray[349] = 12'h369;
iconPixArray[350] = 12'h 11;
iconPixArray[351] = 12'h 00;
iconPixArray[352] = 12'h 00;
iconPixArray[353] = 12'h 00;
iconPixArray[354] = 12'h 00;
iconPixArray[355] = 12'h100;
iconPixArray[356] = 12'h200;
iconPixArray[357] = 12'h100;
iconPixArray[358] = 12'h100;
iconPixArray[359] = 12'h48D;
iconPixArray[360] = 12'h47B;
iconPixArray[361] = 12'h468;
iconPixArray[362] = 12'hBBB;
iconPixArray[363] = 12'hBCC;
iconPixArray[364] = 12'h468;
iconPixArray[365] = 12'h 11;
iconPixArray[366] = 12'h 00;
iconPixArray[367] = 12'h 00;
iconPixArray[368] = 12'h 00;
iconPixArray[369] = 12'h 00;
iconPixArray[370] = 12'h100;
iconPixArray[371] = 12'h600;
iconPixArray[372] = 12'hE00;
iconPixArray[373] = 12'h300;
iconPixArray[374] = 12'h369;
iconPixArray[375] = 12'h677;
iconPixArray[376] = 12'hCCC;
iconPixArray[377] = 12'h457;
iconPixArray[378] = 12'h47A;
iconPixArray[379] = 12'h47A;
iconPixArray[380] = 12'h124;
iconPixArray[381] = 12'h 00;
iconPixArray[382] = 12'h 00;
iconPixArray[383] = 12'h 00;
iconPixArray[384] = 12'h 00;
iconPixArray[385] = 12'h 00;
iconPixArray[386] = 12'h200;
iconPixArray[387] = 12'hE00;
iconPixArray[388] = 12'h700;
iconPixArray[389] = 12'h234;
iconPixArray[390] = 12'h47A;
iconPixArray[391] = 12'hDDD;
iconPixArray[392] = 12'hFFF;
iconPixArray[393] = 12'h788;
iconPixArray[394] = 12'h49E;
iconPixArray[395] = 12'h135;
iconPixArray[396] = 12'h 01;
iconPixArray[397] = 12'h 00;
iconPixArray[398] = 12'h 00;
iconPixArray[399] = 12'h 00;
iconPixArray[400] = 12'h 00;
iconPixArray[401] = 12'h100;
iconPixArray[402] = 12'h900;
iconPixArray[403] = 12'hB00;
iconPixArray[404] = 12'h101;
iconPixArray[405] = 12'h59E;
iconPixArray[406] = 12'h49E;
iconPixArray[407] = 12'h467;
iconPixArray[408] = 12'h788;
iconPixArray[409] = 12'h468;
iconPixArray[410] = 12'h135;
iconPixArray[411] = 12'h 11;
iconPixArray[412] = 12'h 00;
iconPixArray[413] = 12'h 00;
iconPixArray[414] = 12'h 00;
iconPixArray[415] = 12'h 00;
iconPixArray[416] = 12'h 00;
iconPixArray[417] = 12'h 00;
iconPixArray[418] = 12'h100;
iconPixArray[419] = 12'h100;
iconPixArray[420] = 12'h36A;
iconPixArray[421] = 12'h5AF;
iconPixArray[422] = 12'h5AF;
iconPixArray[423] = 12'h5AF;
iconPixArray[424] = 12'h48C;
iconPixArray[425] = 12'h100;
iconPixArray[426] = 12'h100;
iconPixArray[427] = 12'h 00;
iconPixArray[428] = 12'h 00;
iconPixArray[429] = 12'h 00;
iconPixArray[430] = 12'h 00;
iconPixArray[431] = 12'h 00;
iconPixArray[432] = 12'h 00;
iconPixArray[433] = 12'h 00;
iconPixArray[434] = 12'h 00;
iconPixArray[435] = 12'h 00;
iconPixArray[436] = 12'h 01;
iconPixArray[437] = 12'h47B;
iconPixArray[438] = 12'h5AF;
iconPixArray[439] = 12'h36A;
iconPixArray[440] = 12'h100;
iconPixArray[441] = 12'hA00;
iconPixArray[442] = 12'h100;
iconPixArray[443] = 12'h 00;
iconPixArray[444] = 12'h 00;
iconPixArray[445] = 12'h 00;
iconPixArray[446] = 12'h 00;
iconPixArray[447] = 12'h 00;
iconPixArray[448] = 12'h 00;
iconPixArray[449] = 12'h 00;
iconPixArray[450] = 12'h 00;
iconPixArray[451] = 12'h 00;
iconPixArray[452] = 12'h 00;
iconPixArray[453] = 12'h 11;
iconPixArray[454] = 12'h235;
iconPixArray[455] = 12'h200;
iconPixArray[456] = 12'hD00;
iconPixArray[457] = 12'hC00;
iconPixArray[458] = 12'h100;
iconPixArray[459] = 12'h 00;
iconPixArray[460] = 12'h 00;
iconPixArray[461] = 12'h 00;
iconPixArray[462] = 12'h 00;
iconPixArray[463] = 12'h 00;
iconPixArray[464] = 12'h 00;
iconPixArray[465] = 12'h 00;
iconPixArray[466] = 12'h 00;
iconPixArray[467] = 12'h 00;
iconPixArray[468] = 12'h 00;
iconPixArray[469] = 12'h 00;
iconPixArray[470] = 12'h100;
iconPixArray[471] = 12'hE00;
iconPixArray[472] = 12'hC00;
iconPixArray[473] = 12'h100;
iconPixArray[474] = 12'h 00;
iconPixArray[475] = 12'h 00;
iconPixArray[476] = 12'h 00;
iconPixArray[477] = 12'h 00;
iconPixArray[478] = 12'h 00;
iconPixArray[479] = 12'h 00;
iconPixArray[480] = 12'h 00;
iconPixArray[481] = 12'h 00;
iconPixArray[482] = 12'h 00;
iconPixArray[483] = 12'h 00;
iconPixArray[484] = 12'h 00;
iconPixArray[485] = 12'h 00;
iconPixArray[486] = 12'h100;
iconPixArray[487] = 12'h300;
iconPixArray[488] = 12'h100;
iconPixArray[489] = 12'h 00;
iconPixArray[490] = 12'h 00;
iconPixArray[491] = 12'h 00;
iconPixArray[492] = 12'h 00;
iconPixArray[493] = 12'h 00;
iconPixArray[494] = 12'h 00;
iconPixArray[495] = 12'h 00;
iconPixArray[496] = 12'hFFF;
iconPixArray[497] = 12'hFFF;
iconPixArray[498] = 12'hFFF;
iconPixArray[499] = 12'hFFF;
iconPixArray[500] = 12'hFFF;
iconPixArray[501] = 12'hFFF;
iconPixArray[502] = 12'hFFF;
iconPixArray[503] = 12'hFFF;
iconPixArray[504] = 12'hFFF;
iconPixArray[505] = 12'hFFF;
iconPixArray[506] = 12'hFFF;
iconPixArray[507] = 12'hFFF;
iconPixArray[508] = 12'hFFF;
iconPixArray[509] = 12'hFFF;
iconPixArray[510] = 12'hFFF;
iconPixArray[511] = 12'hFFF;
iconPixArray[0] = 12'h 00;
iconPixArray[1] = 12'h 00;
iconPixArray[2] = 12'h 00;
iconPixArray[3] = 12'h 00;
iconPixArray[4] = 12'h 00;
iconPixArray[5] = 12'h 00;
iconPixArray[6] = 12'h 00;
iconPixArray[7] = 12'h 00;
iconPixArray[8] = 12'h 00;
iconPixArray[9] = 12'h 00;
iconPixArray[10] = 12'h 00;
iconPixArray[11] = 12'h 00;
iconPixArray[12] = 12'h 00;
iconPixArray[13] = 12'h 00;
iconPixArray[14] = 12'h 00;
iconPixArray[15] = 12'h 00;
iconPixArray[16] = 12'h 00;
iconPixArray[17] = 12'h 00;
iconPixArray[18] = 12'h 00;
iconPixArray[19] = 12'h 00;
iconPixArray[20] = 12'h 00;
iconPixArray[21] = 12'h 00;
iconPixArray[22] = 12'h 00;
iconPixArray[23] = 12'h 00;
iconPixArray[24] = 12'h 00;
iconPixArray[25] = 12'h 00;
iconPixArray[26] = 12'h 00;
iconPixArray[27] = 12'h 00;
iconPixArray[28] = 12'h 11;
iconPixArray[29] = 12'h 11;
iconPixArray[30] = 12'h 11;
iconPixArray[31] = 12'h 01;
iconPixArray[32] = 12'h 00;
iconPixArray[33] = 12'h 00;
iconPixArray[34] = 12'h 00;
iconPixArray[35] = 12'h 00;
iconPixArray[36] = 12'h 00;
iconPixArray[37] = 12'h 00;
iconPixArray[38] = 12'h 00;
iconPixArray[39] = 12'h 00;
iconPixArray[40] = 12'h 00;
iconPixArray[41] = 12'h 00;
iconPixArray[42] = 12'h 11;
iconPixArray[43] = 12'h124;
iconPixArray[44] = 12'h37A;
iconPixArray[45] = 12'h59E;
iconPixArray[46] = 12'h369;
iconPixArray[47] = 12'h 00;
iconPixArray[48] = 12'h 00;
iconPixArray[49] = 12'h 00;
iconPixArray[50] = 12'h 00;
iconPixArray[51] = 12'h 00;
iconPixArray[52] = 12'h 00;
iconPixArray[53] = 12'h 00;
iconPixArray[54] = 12'h 00;
iconPixArray[55] = 12'h 00;
iconPixArray[56] = 12'h 00;
iconPixArray[57] = 12'h 12;
iconPixArray[58] = 12'h47B;
iconPixArray[59] = 12'h5AF;
iconPixArray[60] = 12'h5AF;
iconPixArray[61] = 12'h5AF;
iconPixArray[62] = 12'h135;
iconPixArray[63] = 12'h 00;
iconPixArray[64] = 12'h 00;
iconPixArray[65] = 12'h 00;
iconPixArray[66] = 12'h 00;
iconPixArray[67] = 12'h 00;
iconPixArray[68] = 12'h 00;
iconPixArray[69] = 12'h 00;
iconPixArray[70] = 12'h 00;
iconPixArray[71] = 12'h 01;
iconPixArray[72] = 12'h123;
iconPixArray[73] = 12'h47B;
iconPixArray[74] = 12'h567;
iconPixArray[75] = 12'h677;
iconPixArray[76] = 12'h47B;
iconPixArray[77] = 12'h59E;
iconPixArray[78] = 12'h 11;
iconPixArray[79] = 12'h 00;
iconPixArray[80] = 12'h 00;
iconPixArray[81] = 12'h 00;
iconPixArray[82] = 12'h 00;
iconPixArray[83] = 12'h 00;
iconPixArray[84] = 12'h 00;
iconPixArray[85] = 12'h 00;
iconPixArray[86] = 12'h 01;
iconPixArray[87] = 12'h123;
iconPixArray[88] = 12'h49E;
iconPixArray[89] = 12'h468;
iconPixArray[90] = 12'hFFF;
iconPixArray[91] = 12'hFFF;
iconPixArray[92] = 12'h568;
iconPixArray[93] = 12'h369;
iconPixArray[94] = 12'h 11;
iconPixArray[95] = 12'h 00;
iconPixArray[96] = 12'h 00;
iconPixArray[97] = 12'h 00;
iconPixArray[98] = 12'h 00;
iconPixArray[99] = 12'h100;
iconPixArray[100] = 12'h200;
iconPixArray[101] = 12'h100;
iconPixArray[102] = 12'h100;
iconPixArray[103] = 12'h48D;
iconPixArray[104] = 12'h47B;
iconPixArray[105] = 12'h468;
iconPixArray[106] = 12'hBBB;
iconPixArray[107] = 12'hBCC;
iconPixArray[108] = 12'h468;
iconPixArray[109] = 12'h 11;
iconPixArray[110] = 12'h 00;
iconPixArray[111] = 12'h 00;
iconPixArray[112] = 12'h 00;
iconPixArray[113] = 12'h 00;
iconPixArray[114] = 12'h100;
iconPixArray[115] = 12'h600;
iconPixArray[116] = 12'hE00;
iconPixArray[117] = 12'h300;
iconPixArray[118] = 12'h369;
iconPixArray[119] = 12'h677;
iconPixArray[120] = 12'hCCC;
iconPixArray[121] = 12'h457;
iconPixArray[122] = 12'h47A;
iconPixArray[123] = 12'h47A;
iconPixArray[124] = 12'h124;
iconPixArray[125] = 12'h 00;
iconPixArray[126] = 12'h 00;
iconPixArray[127] = 12'h 00;
iconPixArray[128] = 12'h 00;
iconPixArray[129] = 12'h 00;
iconPixArray[130] = 12'h200;
iconPixArray[131] = 12'hE00;
iconPixArray[132] = 12'h700;
iconPixArray[133] = 12'h234;
iconPixArray[134] = 12'h47A;
iconPixArray[135] = 12'hDDD;
iconPixArray[136] = 12'hFFF;
iconPixArray[137] = 12'h788;
iconPixArray[138] = 12'h49E;
iconPixArray[139] = 12'h135;
iconPixArray[140] = 12'h 01;
iconPixArray[141] = 12'h 00;
iconPixArray[142] = 12'h 00;
iconPixArray[143] = 12'h 00;
iconPixArray[144] = 12'h 00;
iconPixArray[145] = 12'h100;
iconPixArray[146] = 12'h900;
iconPixArray[147] = 12'hB00;
iconPixArray[148] = 12'h101;
iconPixArray[149] = 12'h59E;
iconPixArray[150] = 12'h49E;
iconPixArray[151] = 12'h467;
iconPixArray[152] = 12'h788;
iconPixArray[153] = 12'h468;
iconPixArray[154] = 12'h135;
iconPixArray[155] = 12'h 11;
iconPixArray[156] = 12'h 00;
iconPixArray[157] = 12'h 00;
iconPixArray[158] = 12'h 00;
iconPixArray[159] = 12'h 00;
iconPixArray[160] = 12'h 00;
iconPixArray[161] = 12'h 00;
iconPixArray[162] = 12'h100;
iconPixArray[163] = 12'h100;
iconPixArray[164] = 12'h36A;
iconPixArray[165] = 12'h5AF;
iconPixArray[166] = 12'h5AF;
iconPixArray[167] = 12'h5AF;
iconPixArray[168] = 12'h48C;
iconPixArray[169] = 12'h100;
iconPixArray[170] = 12'h100;
iconPixArray[171] = 12'h 00;
iconPixArray[172] = 12'h 00;
iconPixArray[173] = 12'h 00;
iconPixArray[174] = 12'h 00;
iconPixArray[175] = 12'h 00;
iconPixArray[176] = 12'h 00;
iconPixArray[177] = 12'h 00;
iconPixArray[178] = 12'h 00;
iconPixArray[179] = 12'h 00;
iconPixArray[180] = 12'h 01;
iconPixArray[181] = 12'h47B;
iconPixArray[182] = 12'h5AF;
iconPixArray[183] = 12'h36A;
iconPixArray[184] = 12'h100;
iconPixArray[185] = 12'hA00;
iconPixArray[186] = 12'h100;
iconPixArray[187] = 12'h 00;
iconPixArray[188] = 12'h 00;
iconPixArray[189] = 12'h 00;
iconPixArray[190] = 12'h 00;
iconPixArray[191] = 12'h 00;
iconPixArray[192] = 12'h 00;
iconPixArray[193] = 12'h 00;
iconPixArray[194] = 12'h 00;
iconPixArray[195] = 12'h 00;
iconPixArray[196] = 12'h 00;
iconPixArray[197] = 12'h 11;
iconPixArray[198] = 12'h235;
iconPixArray[199] = 12'h200;
iconPixArray[200] = 12'hD00;
iconPixArray[201] = 12'hC00;
iconPixArray[202] = 12'h100;
iconPixArray[203] = 12'h 00;
iconPixArray[204] = 12'h 00;
iconPixArray[205] = 12'h 00;
iconPixArray[206] = 12'h 00;
iconPixArray[207] = 12'h 00;
iconPixArray[208] = 12'h 00;
iconPixArray[209] = 12'h 00;
iconPixArray[210] = 12'h 00;
iconPixArray[211] = 12'h 00;
iconPixArray[212] = 12'h 00;
iconPixArray[213] = 12'h 00;
iconPixArray[214] = 12'h100;
iconPixArray[215] = 12'hE00;
iconPixArray[216] = 12'hC00;
iconPixArray[217] = 12'h100;
iconPixArray[218] = 12'h 00;
iconPixArray[219] = 12'h 00;
iconPixArray[220] = 12'h 00;
iconPixArray[221] = 12'h 00;
iconPixArray[222] = 12'h 00;
iconPixArray[223] = 12'h 00;
iconPixArray[224] = 12'h 00;
iconPixArray[225] = 12'h 00;
iconPixArray[226] = 12'h 00;
iconPixArray[227] = 12'h 00;
iconPixArray[228] = 12'h 00;
iconPixArray[229] = 12'h 00;
iconPixArray[230] = 12'h100;
iconPixArray[231] = 12'h300;
iconPixArray[232] = 12'h100;
iconPixArray[233] = 12'h 00;
iconPixArray[234] = 12'h 00;
iconPixArray[235] = 12'h 00;
iconPixArray[236] = 12'h 00;
iconPixArray[237] = 12'h 00;
iconPixArray[238] = 12'h 00;
iconPixArray[239] = 12'h 00;
iconPixArray[240] = 12'hFFF;
iconPixArray[241] = 12'hFFF;
iconPixArray[242] = 12'hFFF;
iconPixArray[243] = 12'hFFF;
iconPixArray[244] = 12'hFFF;
iconPixArray[245] = 12'hFFF;
iconPixArray[246] = 12'hFFF;
iconPixArray[247] = 12'hFFF;
iconPixArray[248] = 12'hFFF;
iconPixArray[249] = 12'hFFF;
iconPixArray[250] = 12'hFFF;
iconPixArray[251] = 12'hFFF;
iconPixArray[252] = 12'hFFF;
iconPixArray[253] = 12'hFFF;
iconPixArray[254] = 12'hFFF;
iconPixArray[255] = 12'hFFF;



end
endmodule 
